magic
tech scmos
timestamp 1598461406
<< nwell >>
rect 46 15 64 36
rect 76 15 94 36
rect 103 15 121 34
rect 130 -10 155 2
<< polysilicon >>
rect 54 26 56 28
rect 84 26 86 28
rect 111 26 113 28
rect 138 27 140 29
rect 54 9 56 16
rect 55 5 56 9
rect 84 6 86 16
rect 111 6 113 16
rect 138 14 140 22
rect 139 10 140 14
rect 54 -2 56 5
rect 85 2 86 6
rect 112 2 113 6
rect 54 -9 56 -7
rect 84 -8 86 2
rect 111 -2 113 2
rect 138 1 140 10
rect 111 -9 113 -7
rect 138 -11 140 -9
rect 84 -15 86 -13
<< ndiffusion >>
rect 131 26 138 27
rect 131 22 132 26
rect 136 22 138 26
rect 140 23 142 27
rect 146 23 147 27
rect 140 22 147 23
rect 47 -6 48 -2
rect 52 -6 54 -2
rect 47 -7 54 -6
rect 56 -6 58 -2
rect 62 -6 63 -2
rect 56 -7 63 -6
rect 104 -6 105 -2
rect 109 -6 111 -2
rect 104 -7 111 -6
rect 113 -6 115 -2
rect 119 -6 120 -2
rect 113 -7 120 -6
rect 77 -12 78 -8
rect 82 -12 84 -8
rect 77 -13 84 -12
rect 86 -12 88 -8
rect 92 -12 93 -8
rect 86 -13 93 -12
<< pdiffusion >>
rect 47 23 54 26
rect 47 19 48 23
rect 52 19 54 23
rect 47 16 54 19
rect 56 23 63 26
rect 56 19 58 23
rect 62 19 63 23
rect 56 16 63 19
rect 77 23 84 26
rect 77 19 78 23
rect 82 19 84 23
rect 77 16 84 19
rect 86 23 93 26
rect 86 19 88 23
rect 92 19 93 23
rect 86 16 93 19
rect 104 23 111 26
rect 104 19 105 23
rect 109 19 111 23
rect 104 16 111 19
rect 113 23 120 26
rect 113 19 115 23
rect 119 19 120 23
rect 113 16 120 19
rect 131 -2 138 1
rect 131 -6 132 -2
rect 136 -6 138 -2
rect 131 -9 138 -6
rect 140 -2 147 1
rect 140 -6 142 -2
rect 146 -6 147 -2
rect 140 -9 147 -6
<< metal1 >>
rect 52 30 56 34
rect 60 30 78 34
rect 82 30 86 34
rect 90 30 92 34
rect 101 30 105 34
rect 109 30 146 34
rect 48 23 52 30
rect 78 23 82 30
rect 105 23 109 30
rect 142 27 146 30
rect 49 5 51 9
rect 58 6 62 19
rect 88 13 92 19
rect 92 9 100 13
rect 115 6 119 19
rect 132 20 136 22
rect 132 17 146 20
rect 126 10 135 13
rect 126 9 139 10
rect 142 11 146 17
rect 142 8 160 11
rect 142 6 146 8
rect 58 2 81 6
rect 85 2 108 6
rect 115 2 146 6
rect 58 -2 62 2
rect 115 -2 119 2
rect 142 -2 146 2
rect 151 2 155 8
rect 48 -18 52 -6
rect 88 -8 92 -5
rect 105 -11 109 -6
rect 132 -11 136 -6
rect 78 -18 82 -12
rect 101 -15 136 -11
rect 52 -22 56 -18
rect 60 -22 78 -18
rect 82 -22 86 -18
rect 90 -22 91 -18
<< metal2 >>
rect 104 9 122 13
rect 88 -1 92 9
<< ntransistor >>
rect 138 22 140 27
rect 54 -7 56 -2
rect 111 -7 113 -2
rect 84 -13 86 -8
<< ptransistor >>
rect 54 16 56 26
rect 84 16 86 26
rect 111 16 113 26
rect 138 -9 140 1
<< polycontact >>
rect 51 5 55 9
rect 135 10 139 14
rect 81 2 85 6
rect 108 2 112 6
<< ndcontact >>
rect 132 22 136 26
rect 142 23 146 27
rect 48 -6 52 -2
rect 58 -6 62 -2
rect 105 -6 109 -2
rect 115 -6 119 -2
rect 78 -12 82 -8
rect 88 -12 92 -8
<< pdcontact >>
rect 48 19 52 23
rect 58 19 62 23
rect 78 19 82 23
rect 88 19 92 23
rect 105 19 109 23
rect 115 19 119 23
rect 132 -6 136 -2
rect 142 -6 146 -2
<< m2contact >>
rect 88 9 92 13
rect 100 9 104 13
rect 122 9 126 13
rect 88 -5 92 -1
<< psubstratepcontact >>
rect 48 -22 52 -18
rect 56 -22 60 -18
rect 78 -22 82 -18
rect 86 -22 90 -18
<< nsubstratencontact >>
rect 48 30 52 34
rect 56 30 60 34
rect 78 30 82 34
rect 86 30 90 34
rect 105 30 109 34
rect 151 -2 155 2
<< labels >>
rlabel metal1 49 5 49 9 3 digital_input
rlabel metal1 101 30 101 34 5 V_in1
rlabel metal1 101 -15 101 -11 1 V_in2
rlabel metal1 64 4 64 4 1 dig_inv
rlabel metal1 84 -20 84 -20 1 gnd!
rlabel metal1 54 -20 54 -20 1 gnd!
rlabel metal1 97 10 97 10 1 dig_inv_inv
rlabel metal1 160 8 160 11 7 V_out
rlabel metal1 62 32 62 32 5 v1
<< end >>
