* SPICE3 file created from 8BitDac.ext - technology: scmos


.model polyResistor R ( TC1=0 TC2=0 RSH=7.7 DEFW=1.E-7 NARROW=0.0 TNOM=27)

.model pfet PMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=4.1589E17 VTH0=-0.3938813 K1=0.5479015 K2=0.0360586 K3=0.0993095 K3B=5.7086622 W0=1E-6 NLX=1.313191E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=0.4911363 DVT1=0.2227356 DVT2=0.1 U0=115.6852975 UA=1.505832E-9 UB=1E-21 UC=-1E-10 VSAT=1.329694E5 A0=1.7590478 AGS=0.3641621 B0=3.427126E-7 B1=1.062928E-6 KETA=0.0134667 A1=0.6859506 A2=0.3506788 RDSW=168.5705677 PRWG=0.5 PRWB=-0.4987371 WR=1 WINT=0 LINT=3.028832E-8 XL=0 XW=-1E-8 DWG=-2.349633E-8 DWB=-7.152486E-9 VOFF=-0.0994037 NFACTOR=1.9424315 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=0.0608072 ETAB=-0.0426148 DSUB=0.7343015 PCLM=3.2579974 PDIBLC1=7.229527E-6 PDIBLC2=0.025389 PDIBLCB=-1E-3 DROUT=0 PSCBE1=1.454878E10 PSCBE2=4.202027E-9 PVAG=15 DELTA=0.01 RSH=7.8 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=6.32E-10 CGSO=6.32E-10 CGBO=1E-12 CJ=1.172138E-3 PB=0.8421173 MJ=0.4109788 CJSW=2.242609E-10 PBSW=0.8 MJSW=0.3752089 CJSWG=4.22E-10 PBSWG=0.8 MJSWG=0.3752089 CF=0 PVTH0=1.888482E-3 PRDSW=11.5315407 PK2=1.559399E-3 WKETA=0.0319301 LKETA=2.955547E-3 PU0=-1.1105313 PUA=-4.62102E-11 PUB=1E-21 PVSAT=50 PETA0=1E-4 PKETA=-4.346368E-3)

.model nfet NMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=2.3549E17 VTH0=0.3823463 K1=0.5810697 K2=4.774618E-3 K3=0.0431669 K3B=1.1498346 W0=1E-7 NLX=1.910552E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=1.2894824 DVT1=0.3622063 DVT2=0.0713729 U0=280.633249 UA=-1.208537E-9 UB=2.158625E-18 UC=5.342807E-11 VSAT=9.366802E4 A0=1.7593146 AGS=0.3939741 B0=-6.413949E-9 B1=-1E-7 KETA=-5.180424E-4 A1=0 A2=1 RDSW=105.5517558 PRWG=0.5 PRWB=-0.1998871 WR=1 WINT=7.904732E-10 LINT=1.571424E-8 XL=0 XW=-1E-8 DWG=1.297221E-9 DWB=1.479041E-9 VOFF=-0.0955434 NFACTOR=2.4358891 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=3.104851E-3 ETAB=-2.512384E-5 DSUB=0.0167075 PCLM=0.8073191 PDIBLC1=0.1666161 PDIBLC2=3.112892E-3 PDIBLCB=-0.1 DROUT=0.7875618 PSCBE1=8E10 PSCBE2=9.213635E-10 PVAG=3.85243E-3 DELTA=0.01 RSH=6.7 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=7.08E-10 CGSO=7.08E-10 CGBO=1E-12 CJ=9.68858E-4 PB=0.8 MJ=0.3864502 CJSW=2.512138E-10 PBSW=0.809286 MJSW=0.1060414 CJSWG=3.3E-10 PBSWG=0.809286 MJSWG=0.1060414 CF=0 PVTH0=-1.192722E-3 PRDSW=-5 PK2=6.450505E-5 WKETA=-4.27294E-4 LKETA=-0.0104078 PU0=6.3268729 PUA=2.226552E-11 PUB=0 PVSAT=969.1480157 PETA0=1E-4 PKETA=-1.049509E-3)





.option scale=0.1u

M1000 7BitDac_1/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=35700 ps=17340
M1001 7BitDac_1/switchNew_0/a_105_21# 7BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1002 7BitDac_1/V_out7 7BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/V_out6 7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1003 7BitDac_1/6BitDac_0/V_out6 7BitDac_1/switchNew_0/a_105_21# 7BitDac_1/V_out7 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1004 7BitDac_1/switchNew_0/a_86_24# D6 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=17850 ps=12240
M1005 7BitDac_1/switchNew_0/a_105_21# 7BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1006 7BitDac_1/V_out7 7BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/V_out6 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1007 7BitDac_1/V_out7 7BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/V_out6 7BitDac_1/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1008 7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1009 7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1010 7BitDac_1/6BitDac_1/V_out6 7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/V_out5 7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1011 7BitDac_1/6BitDac_1/5BitDac_0/V_out5 7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/V_out6 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1012 7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1013 7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1014 7BitDac_1/6BitDac_1/V_out6 7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/V_out5 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1015 7BitDac_1/6BitDac_1/V_out6 7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/V_out5 7BitDac_1/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1016 7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1017 7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1018 7BitDac_1/6BitDac_1/5BitDac_1/V_out5 7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1019 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/V_out5 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1020 7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1021 7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1022 7BitDac_1/6BitDac_1/5BitDac_1/V_out5 7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1023 7BitDac_1/6BitDac_1/5BitDac_1/V_out5 7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 7BitDac_1/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1024 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1025 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1026 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1027 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1028 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1029 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1030 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1031 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1032 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1033 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1034 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1035 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1036 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1037 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1038 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# R_out8 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1039 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# R_out8 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R0 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma R_out8 polyResistor w=2 l=62
M1040 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1041 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1042 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1043 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1044 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1045 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1046 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1047 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1048 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1049 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1050 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1051 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1052 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1053 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1054 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1057 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1058 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1059 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1060 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1061 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1062 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1063 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1064 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1065 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1066 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1067 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1068 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1069 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1070 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1071 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R4 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1072 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1073 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1074 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1075 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1076 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1077 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1078 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1079 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R5 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R6 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R7 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1080 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1081 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1082 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1083 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1084 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1085 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1086 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1089 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1090 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1091 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1092 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1093 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1094 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1095 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1096 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1097 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1098 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1099 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1100 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1101 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1102 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1103 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R8 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M1104 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1105 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1106 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1107 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1108 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1109 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1110 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1111 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R9 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R10 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R11 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1112 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1113 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1114 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1115 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1116 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1117 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1118 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1121 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1122 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1123 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1124 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1125 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1126 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1127 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1128 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1129 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1130 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1131 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1132 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1133 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1134 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1135 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R12 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1136 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1137 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1138 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1139 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1140 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1141 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1142 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1143 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R13 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R14 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R15 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1144 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1145 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1146 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1147 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1148 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1149 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1150 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1151 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1152 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1153 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1154 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1155 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1156 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1157 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1158 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1159 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R16 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M1160 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1161 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1162 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1163 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1164 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1165 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1166 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1167 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R17 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R18 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R19 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1168 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1169 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1170 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1171 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1172 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1173 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1174 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1177 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1178 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1179 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1180 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1181 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1182 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1183 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1184 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1185 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1186 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1187 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1188 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1189 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1190 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1191 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R20 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1192 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1193 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1194 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1195 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1196 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1197 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1198 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1199 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R21 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R22 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R23 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1200 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1201 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1202 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1203 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1204 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1205 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1206 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1209 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1210 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1211 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1212 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1213 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1214 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1215 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1216 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1217 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1218 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1219 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1220 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1221 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1222 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1223 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R24 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M1224 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1225 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1226 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1227 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1228 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1229 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1230 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1231 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R25 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R26 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R27 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1232 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1233 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1234 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1235 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1236 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1237 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1238 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1240 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1241 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1242 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1243 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1244 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1245 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1246 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1247 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1248 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1249 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1250 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1251 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1252 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1253 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1254 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1255 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R28 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1256 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1257 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1258 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1259 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1260 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1261 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1262 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1263 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R29 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R30 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R31 7BitDac_1/6BitDac_1/5BitDac_1/R_in5 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1264 7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1265 7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1266 7BitDac_1/6BitDac_1/5BitDac_0/V_out5 7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1267 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/V_out5 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1268 7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1269 7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1270 7BitDac_1/6BitDac_1/5BitDac_0/V_out5 7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1271 7BitDac_1/6BitDac_1/5BitDac_0/V_out5 7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1272 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1273 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1274 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1275 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1276 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1277 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1278 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1279 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1280 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1281 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1282 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1283 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1284 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1285 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1286 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_1/R_in5 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1287 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_1/R_in5 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R32 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M1288 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1289 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1290 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1291 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1292 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1293 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1294 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1295 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R33 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R34 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R35 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1296 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1297 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1298 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1299 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1300 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1301 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1302 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1303 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1304 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1305 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1306 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1307 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1308 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1309 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1310 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1311 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1312 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1313 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1314 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1315 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1316 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1317 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1318 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1319 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R36 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1320 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1321 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1322 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1323 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1324 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1325 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1326 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1327 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R37 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R38 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R39 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1328 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1329 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1330 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1331 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1332 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1333 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1334 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1335 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1336 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1337 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1338 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1339 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1340 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1341 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1342 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1343 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1344 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1345 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1346 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1347 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1348 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1349 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1350 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1351 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R40 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M1352 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1353 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1354 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1355 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1356 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1357 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1358 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1359 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R41 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R42 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R43 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1360 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1361 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1362 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1363 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1364 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1365 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1366 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1367 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1368 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1369 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1370 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1371 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1372 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1373 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1374 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1375 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1376 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1377 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1378 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1379 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1380 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1381 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1382 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1383 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R44 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1384 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1385 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1386 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1387 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1388 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1389 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1390 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1391 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R45 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R46 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R47 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1392 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1393 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1394 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1395 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1396 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1397 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1398 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1399 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1400 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1401 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1402 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1403 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1404 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1405 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1406 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1407 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R48 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M1408 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1409 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1410 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1411 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1412 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1413 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1414 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1415 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R49 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R50 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R51 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1416 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1417 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1418 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1419 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1420 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1421 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1422 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1423 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1424 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1425 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1426 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1427 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1428 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1429 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1430 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1431 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1432 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1433 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1434 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1435 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1436 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1437 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1438 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1439 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R52 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1440 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1441 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1442 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1443 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1444 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1445 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1446 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1447 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R53 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R54 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R55 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1448 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1449 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1450 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1451 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1452 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1453 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1454 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1455 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1456 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1457 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1458 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1459 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1460 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1461 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1462 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1463 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1464 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1465 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1466 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1467 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1468 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1469 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1470 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1471 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R56 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M1472 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1473 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1474 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1475 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1476 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1477 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1478 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1479 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R57 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R58 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R59 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1480 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1481 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1482 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1483 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1484 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1485 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1486 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1487 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1488 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1489 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1490 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1491 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1492 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1493 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1494 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1495 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1496 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1497 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1498 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1499 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1500 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1501 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1502 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1503 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R60 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1504 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1505 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1506 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1507 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1508 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1509 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1510 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1511 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R61 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R62 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R63 7BitDac_1/6BitDac_1/R_in6 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1512 7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1513 7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1514 7BitDac_1/6BitDac_0/V_out6 7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/V_out5 7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1515 7BitDac_1/6BitDac_0/5BitDac_0/V_out5 7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/V_out6 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1516 7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1517 7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1518 7BitDac_1/6BitDac_0/V_out6 7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/V_out5 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1519 7BitDac_1/6BitDac_0/V_out6 7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/V_out5 7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1520 7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1521 7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1522 7BitDac_1/6BitDac_0/5BitDac_1/V_out5 7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1523 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/V_out5 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1524 7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1525 7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1526 7BitDac_1/6BitDac_0/5BitDac_1/V_out5 7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1527 7BitDac_1/6BitDac_0/5BitDac_1/V_out5 7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 7BitDac_1/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1528 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1529 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1530 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1531 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1532 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1533 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1534 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1535 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1536 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1537 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1538 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1539 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1540 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1541 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1542 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_1/R_in6 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1543 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_1/R_in6 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R64 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_1/R_in6 polyResistor w=2 l=62
M1544 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1545 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1546 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1547 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1548 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1549 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1550 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1551 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R65 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R66 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R67 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1552 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1553 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1554 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1555 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1556 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1557 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1558 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1559 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1560 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1561 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1562 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1563 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1564 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1565 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1566 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1567 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1568 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1569 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1570 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1571 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1572 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1573 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1574 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1575 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R68 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1576 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1577 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1578 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1579 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1580 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1581 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1582 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1583 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R69 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R70 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R71 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1584 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1585 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1586 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1587 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1588 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1589 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1590 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1591 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1592 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1593 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1594 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1595 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1596 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1597 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1598 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1599 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1600 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1601 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1602 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1603 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1604 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1605 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1606 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1607 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R72 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M1608 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1609 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1610 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1611 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1612 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1613 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1614 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1615 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R73 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R74 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R75 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1616 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1617 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1618 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1619 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1620 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1621 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1622 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1623 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1624 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1625 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1626 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1627 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1628 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1629 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1630 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1631 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1632 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1633 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1634 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1635 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1636 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1637 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1638 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1639 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R76 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1640 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1641 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1642 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1643 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1644 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1645 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1646 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1647 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R77 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R78 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R79 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1648 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1649 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1650 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1651 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1652 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1653 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1654 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1655 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1656 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1657 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1658 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1659 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1660 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1661 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1662 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1663 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R80 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M1664 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1665 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1666 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1667 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1668 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1669 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1670 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1671 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R81 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R82 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R83 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1672 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1673 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1674 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1675 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1676 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1677 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1678 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1679 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1680 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1681 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1682 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1683 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1684 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1685 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1686 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1687 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1688 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1689 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1690 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1691 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1692 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1693 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1694 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1695 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R84 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1696 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1697 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1698 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1699 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1700 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1701 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1702 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1703 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R85 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R86 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R87 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1704 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1705 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1706 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1707 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1708 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1709 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1710 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1711 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1712 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1713 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1714 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1715 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1716 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1717 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1718 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1719 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1720 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1721 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1722 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1723 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1724 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1725 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1726 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1727 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R88 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M1728 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1729 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1730 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1731 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1732 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1733 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1734 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1735 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R89 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R90 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R91 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1736 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1737 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1738 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1739 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1740 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1741 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1742 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1743 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1744 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1745 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1746 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1747 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1748 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1749 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1750 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1751 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1752 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1753 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1754 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1755 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1756 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1757 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1758 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1759 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R92 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1760 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1761 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1762 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1763 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1764 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1765 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1766 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1767 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R93 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R94 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R95 7BitDac_1/6BitDac_0/5BitDac_1/R_in5 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1768 7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1769 7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1770 7BitDac_1/6BitDac_0/5BitDac_0/V_out5 7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1771 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/V_out5 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1772 7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1773 7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1774 7BitDac_1/6BitDac_0/5BitDac_0/V_out5 7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1775 7BitDac_1/6BitDac_0/5BitDac_0/V_out5 7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1776 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1777 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1778 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1779 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1780 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1781 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1782 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1783 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1784 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1785 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1786 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1787 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1788 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1789 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1790 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_1/R_in5 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1791 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_1/R_in5 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R96 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M1792 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1793 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1794 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1795 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1796 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1797 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1798 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1799 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R97 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R98 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R99 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1800 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1801 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1802 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1803 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1804 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1805 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1806 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1807 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1808 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1809 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1810 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1811 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1812 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1813 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1814 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1815 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1816 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1817 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1818 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1819 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1820 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1821 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1822 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1823 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R100 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1824 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1825 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1826 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1827 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1828 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1829 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1830 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1831 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R101 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R102 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R103 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1832 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1833 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1834 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1835 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1836 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1837 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1838 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1839 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1840 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1841 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1842 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1843 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1844 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1845 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1846 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1847 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1848 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1849 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1850 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1851 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1852 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1853 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1854 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1855 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R104 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M1856 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1857 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1858 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1859 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1860 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1861 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1862 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1863 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R105 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R106 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R107 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1864 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1865 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1866 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1867 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1868 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1869 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1870 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1871 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1872 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1873 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1874 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1875 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1876 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1877 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1878 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1879 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1880 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1881 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1882 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1883 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1884 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1885 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1886 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1887 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R108 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1888 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1889 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1890 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1891 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1892 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1893 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1894 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1895 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R109 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R110 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R111 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1896 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1897 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1898 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1899 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1900 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1901 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1902 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1903 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1904 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1905 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1906 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1907 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1908 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1909 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1910 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1911 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R112 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M1912 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1913 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1914 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1915 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1916 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1917 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1918 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1919 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R113 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R114 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R115 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1920 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1921 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1922 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1923 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1924 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1925 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1926 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1927 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1928 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1929 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1930 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1931 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1932 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1933 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1934 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1935 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1936 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1937 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1938 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1939 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1940 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1941 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1942 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1943 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R116 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1944 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1945 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1946 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1947 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1948 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1949 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1950 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1951 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R117 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R118 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R119 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1952 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1953 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1954 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1955 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1956 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1957 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1958 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1959 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1960 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1961 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1962 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1963 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1964 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1965 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1966 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1967 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1968 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1969 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1970 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1971 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1972 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1973 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1974 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1975 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R120 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M1976 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1977 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1978 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1979 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1980 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1981 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1982 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1983 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R121 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R122 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R123 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1984 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1985 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1986 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1987 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1988 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1989 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1990 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1991 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1992 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1993 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1994 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1995 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1996 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1997 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1998 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1999 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2000 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2001 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2002 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2003 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2004 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2005 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2006 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2007 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R124 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2008 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2009 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2010 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2011 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2012 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2013 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2014 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2015 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R125 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R126 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R127 7BitDac_1/R_in7 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2016 switchNew_0/a_86_24# D7 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2017 switchNew_0/a_105_21# switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2018 V_out8 switchNew_0/a_86_24# 7BitDac_0/V_out7 7BitDac_0/V_out7 pfet w=10 l=2
+  ad=140 pd=68 as=210 ps=102
M2019 7BitDac_0/V_out7 switchNew_0/a_105_21# V_out8 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=86 ps=64
M2020 switchNew_0/a_86_24# D7 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2021 switchNew_0/a_105_21# switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2022 V_out8 switchNew_0/a_86_24# 7BitDac_1/V_out7 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2023 V_out8 switchNew_0/a_105_21# 7BitDac_1/V_out7 V_out8 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2024 7BitDac_0/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2025 7BitDac_0/switchNew_0/a_105_21# 7BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2026 7BitDac_0/V_out7 7BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/V_out6 7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2027 7BitDac_0/6BitDac_0/V_out6 7BitDac_0/switchNew_0/a_105_21# 7BitDac_0/V_out7 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2028 7BitDac_0/switchNew_0/a_86_24# D6 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2029 7BitDac_0/switchNew_0/a_105_21# 7BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2030 7BitDac_0/V_out7 7BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/V_out6 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2031 7BitDac_0/V_out7 7BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/V_out6 7BitDac_0/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2032 7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2033 7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2034 7BitDac_0/6BitDac_1/V_out6 7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/V_out5 7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2035 7BitDac_0/6BitDac_1/5BitDac_0/V_out5 7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/V_out6 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2036 7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2037 7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2038 7BitDac_0/6BitDac_1/V_out6 7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/V_out5 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2039 7BitDac_0/6BitDac_1/V_out6 7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/V_out5 7BitDac_0/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2040 7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2041 7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2042 7BitDac_0/6BitDac_1/5BitDac_1/V_out5 7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2043 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/V_out5 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2044 7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2045 7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2046 7BitDac_0/6BitDac_1/5BitDac_1/V_out5 7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2047 7BitDac_0/6BitDac_1/5BitDac_1/V_out5 7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 7BitDac_0/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2048 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2049 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2050 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2051 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2052 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2053 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2054 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2055 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2056 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2057 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2058 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2059 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2060 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2061 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2062 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_1/R_in7 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2063 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_1/R_in7 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R128 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_1/R_in7 polyResistor w=2 l=62
M2064 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2065 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2066 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2067 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2068 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2069 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2070 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2071 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R129 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R130 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R131 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2072 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2073 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2074 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2075 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2076 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2077 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2078 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2079 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2080 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2081 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2082 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2083 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2084 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2085 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2086 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2087 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2088 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2089 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2090 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2091 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2092 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2093 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2094 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2095 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R132 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2096 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2097 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2098 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2099 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2100 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2101 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2102 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2103 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R133 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R134 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R135 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2104 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2105 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2106 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2107 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2108 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2109 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2110 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2111 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2112 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2113 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2114 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2115 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2116 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2117 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2118 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2119 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2120 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2121 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2122 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2123 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2124 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2125 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2126 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2127 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R136 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M2128 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2129 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2130 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2131 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2132 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2133 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2134 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2135 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R137 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R138 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R139 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2136 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2137 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2138 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2139 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2140 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2141 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2142 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2143 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2144 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2145 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2146 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2147 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2148 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2149 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2150 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2151 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2152 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2153 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2154 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2155 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2156 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2157 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2158 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2159 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R140 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2160 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2161 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2162 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2163 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2164 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2165 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2166 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2167 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R141 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R142 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R143 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2168 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2169 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2170 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2171 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2172 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2173 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2174 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2175 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2176 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2177 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2178 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2179 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2180 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2181 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2182 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2183 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R144 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M2184 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2185 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2186 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2187 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2188 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2189 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2190 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2191 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R145 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R146 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R147 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2192 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2193 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2194 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2195 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2196 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2197 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2198 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2199 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2200 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2201 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2202 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2203 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2204 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2205 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2206 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2207 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2208 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2209 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2210 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2211 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2212 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2213 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2214 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2215 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R148 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2216 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2217 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2218 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2219 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2220 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2221 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2222 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2223 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R149 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R150 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R151 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2224 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2225 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2226 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2227 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2228 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2229 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2230 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2231 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2232 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2233 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2234 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2235 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2236 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2237 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2238 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2239 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2240 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2241 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2242 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2243 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2244 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2245 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2246 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2247 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R152 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M2248 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2249 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2250 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2251 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2252 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2253 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2254 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2255 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R153 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R154 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R155 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2256 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2257 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2258 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2259 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2260 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2261 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2262 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2263 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2264 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2265 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2266 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2267 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2268 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2269 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2270 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2271 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2272 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2273 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2274 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2275 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2276 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2277 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2278 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2279 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R156 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2280 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2281 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2282 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2283 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2284 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2285 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2286 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2287 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R157 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R158 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R159 7BitDac_0/6BitDac_1/5BitDac_1/R_in5 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2288 7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2289 7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2290 7BitDac_0/6BitDac_1/5BitDac_0/V_out5 7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2291 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/V_out5 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2292 7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2293 7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2294 7BitDac_0/6BitDac_1/5BitDac_0/V_out5 7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2295 7BitDac_0/6BitDac_1/5BitDac_0/V_out5 7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2296 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2297 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2298 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2299 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2300 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2301 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2302 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2303 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2304 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2305 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2306 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2307 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2308 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2309 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2310 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_1/R_in5 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2311 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_1/R_in5 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R160 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M2312 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2313 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2314 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2315 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2316 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2317 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2318 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2319 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R161 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R162 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R163 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2320 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2321 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2322 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2323 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2324 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2325 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2326 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2327 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2328 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2329 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2330 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2331 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2332 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2333 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2334 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2335 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2336 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2337 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2338 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2339 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2340 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2341 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2342 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2343 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R164 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2344 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2345 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2346 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2347 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2348 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2349 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2350 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2351 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R165 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R166 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R167 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2352 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2353 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2354 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2355 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2356 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2357 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2358 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2359 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2360 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2361 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2362 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2363 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2364 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2365 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2366 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2367 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2368 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2369 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2370 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2371 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2372 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2373 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2374 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2375 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R168 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M2376 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2377 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2378 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2379 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2380 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2381 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2382 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2383 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R169 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R170 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R171 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2384 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2385 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2386 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2387 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2388 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2389 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2390 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2391 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2392 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2393 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2394 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2395 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2396 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2397 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2398 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2399 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2400 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2401 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2402 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2403 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2404 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2405 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2406 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2407 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R172 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2408 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2409 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2410 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2411 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2412 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2413 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2414 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2415 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R173 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R174 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R175 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2416 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2417 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2418 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2419 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2420 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2421 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2422 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2423 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2424 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2425 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2426 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2427 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2428 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2429 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2430 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2431 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R176 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M2432 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2433 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2434 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2435 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2436 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2437 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2438 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2439 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R177 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R178 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R179 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2440 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2441 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2442 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2443 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2444 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2445 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2446 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2447 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2448 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2449 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2450 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2451 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2452 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2453 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2454 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2455 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2456 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2457 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2458 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2459 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2460 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2461 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2462 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2463 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R180 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2464 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2465 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2466 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2467 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2468 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2469 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2470 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2471 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R181 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R182 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R183 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2472 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2473 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2474 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2475 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2476 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2477 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2478 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2479 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2480 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2481 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2482 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2483 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2484 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2485 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2486 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2487 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2488 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2489 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2490 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2491 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2492 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2493 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2494 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2495 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R184 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M2496 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2497 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2498 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2499 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2500 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2501 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2502 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2503 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R185 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R186 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R187 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2504 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2505 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2506 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2507 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2508 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2509 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2510 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2511 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2512 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2513 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2514 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2515 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2516 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2517 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2518 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2519 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2520 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2521 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2522 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2523 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2524 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2525 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2526 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2527 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R188 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2528 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2529 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2530 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2531 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2532 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2533 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2534 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2535 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R189 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R190 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R191 7BitDac_0/6BitDac_1/R_in6 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2536 7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2537 7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2538 7BitDac_0/6BitDac_0/V_out6 7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/V_out5 7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2539 7BitDac_0/6BitDac_0/5BitDac_0/V_out5 7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/V_out6 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2540 7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2541 7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2542 7BitDac_0/6BitDac_0/V_out6 7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/V_out5 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2543 7BitDac_0/6BitDac_0/V_out6 7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/V_out5 7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2544 7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2545 7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2546 7BitDac_0/6BitDac_0/5BitDac_1/V_out5 7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2547 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/V_out5 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2548 7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2549 7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2550 7BitDac_0/6BitDac_0/5BitDac_1/V_out5 7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2551 7BitDac_0/6BitDac_0/5BitDac_1/V_out5 7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 7BitDac_0/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2552 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2553 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2554 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2555 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2556 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2557 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2558 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2559 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2560 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2561 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2562 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2563 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2564 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2565 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2566 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_1/R_in6 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2567 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_1/R_in6 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R192 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_1/R_in6 polyResistor w=2 l=62
M2568 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2569 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2570 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2571 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2572 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2573 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2574 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2575 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R193 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R194 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R195 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2576 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2577 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2578 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2579 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2580 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2581 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2582 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2583 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2584 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2585 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2586 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2587 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2588 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2589 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2590 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2591 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2592 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2593 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2594 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2595 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2596 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2597 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2598 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2599 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R196 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2600 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2601 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2602 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2603 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2604 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2605 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2606 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2607 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R197 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R198 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R199 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2608 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2609 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2610 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2611 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2612 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2613 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2614 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2615 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2616 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2617 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2618 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2619 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2620 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2621 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2622 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2623 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2624 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2625 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2626 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2627 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2628 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2629 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2630 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2631 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R200 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M2632 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2633 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2634 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2635 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2636 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2637 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2638 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2639 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R201 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R202 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R203 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2640 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2641 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2642 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2643 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2644 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2645 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2646 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2647 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2648 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2649 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2650 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2651 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2652 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2653 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2654 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2655 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2656 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2657 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2658 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2659 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2660 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2661 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2662 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2663 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R204 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2664 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2665 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2666 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2667 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2668 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2669 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2670 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2671 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R205 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R206 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R207 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2672 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2673 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2674 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2675 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2676 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2677 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2678 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2679 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2680 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2681 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2682 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2683 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2684 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2685 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2686 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2687 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R208 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M2688 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2689 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2690 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2691 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2692 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2693 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2694 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2695 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R209 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R210 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R211 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2696 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2697 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2698 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2699 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2700 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2701 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2702 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2703 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2704 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2705 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2706 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2707 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2708 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2709 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2710 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2711 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2712 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2713 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2714 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2715 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2716 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2717 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2718 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2719 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R212 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2720 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2721 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2722 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2723 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2724 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2725 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2726 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2727 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R213 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R214 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R215 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2728 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2729 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2730 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2731 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2732 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2733 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2734 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2735 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2736 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2737 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2738 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2739 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2740 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2741 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2742 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2743 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2744 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2745 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2746 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2747 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2748 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2749 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2750 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2751 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R216 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M2752 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2753 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2754 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2755 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2756 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2757 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2758 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2759 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R217 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R218 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R219 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2760 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2761 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2762 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2763 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2764 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2765 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2766 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2767 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2768 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2769 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2770 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2771 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2772 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2773 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2774 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2775 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2776 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2777 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2778 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2779 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2780 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2781 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2782 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2783 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R220 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2784 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2785 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2786 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2787 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2788 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2789 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2790 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2791 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R221 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R222 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R223 7BitDac_0/6BitDac_0/5BitDac_1/R_in5 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2792 7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2793 7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2794 7BitDac_0/6BitDac_0/5BitDac_0/V_out5 7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2795 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/V_out5 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2796 7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2797 7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2798 7BitDac_0/6BitDac_0/5BitDac_0/V_out5 7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2799 7BitDac_0/6BitDac_0/5BitDac_0/V_out5 7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2800 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2801 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2802 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2803 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2804 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2805 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2806 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2807 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2808 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2809 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2810 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2811 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2812 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2813 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2814 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_1/R_in5 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2815 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_1/R_in5 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R224 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M2816 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2817 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2818 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2819 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2820 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2821 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2822 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2823 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R225 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R226 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R227 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2824 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2825 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2826 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2827 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2828 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2829 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2830 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2831 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2832 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2833 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2834 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2835 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2836 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2837 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2838 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2839 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2840 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2841 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2842 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2843 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2844 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2845 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2846 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2847 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R228 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2848 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2849 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2850 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2851 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2852 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2853 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2854 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2855 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R229 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R230 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R231 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2856 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2857 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2858 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2859 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2860 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2861 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2862 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2863 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2864 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2865 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2866 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2867 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2868 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2869 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2870 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2871 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2872 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2873 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2874 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2875 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2876 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2877 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2878 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2879 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R232 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M2880 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2881 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2882 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2883 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2884 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2885 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2886 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2887 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R233 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R234 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R235 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2888 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2889 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2890 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2891 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2892 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2893 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2894 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2895 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2896 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2897 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2898 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2899 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2900 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2901 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2902 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2903 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2904 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2905 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2906 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2907 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2908 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2909 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2910 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2911 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R236 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2912 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2913 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2914 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2915 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2916 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2917 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2918 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2919 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R237 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R238 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R239 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2920 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2921 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2922 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2923 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2924 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2925 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2926 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2927 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2928 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2929 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2930 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2931 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2932 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2933 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2934 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2935 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R240 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M2936 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2937 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2938 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2939 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2940 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2941 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2942 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2943 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R241 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R242 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R243 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2944 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2945 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2946 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2947 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2948 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2949 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2950 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2951 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2952 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2953 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2954 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2955 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2956 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2957 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2958 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2959 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2960 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2961 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2962 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2963 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2964 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2965 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2966 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2967 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R244 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2968 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2969 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2970 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2971 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2972 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2973 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2974 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2975 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R245 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R246 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R247 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2976 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2977 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2978 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2979 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2980 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2981 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2982 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2983 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2984 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2985 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2986 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2987 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2988 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2989 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2990 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2991 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2992 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2993 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2994 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2995 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2996 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2997 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2998 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2999 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R248 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M3000 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3001 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3002 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3003 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3004 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3005 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3006 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3007 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R249 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R250 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R251 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3008 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3009 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3010 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3011 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3012 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3013 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3014 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3015 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3016 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3017 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3018 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3019 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3020 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3021 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3022 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3023 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3024 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3025 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3026 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3027 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3028 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3029 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3030 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3031 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R252 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3032 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3033 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3034 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3035 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# m6_733_n10# nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3036 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3037 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# m6_733_n10# m6_733_n10# nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3038 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta m6_733_n10# nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3039 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R253 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R254 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R255 R_in8 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
C0 D2 D1 58.15fF
C1 VA D1 30.50fF
C2 D0 VA 10.36fF
C3 D6 7BitDac_0/6BitDac_0/V_out6 5.31fF
C4 D3 D1 11.09fF
C5 D2 VA 11.38fF
C6 D6 7BitDac_1/6BitDac_0/V_out6 5.31fF
C7 VA D3 15.73fF
C8 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C9 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C10 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C11 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C12 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 m6_733_n10# 2.39fF
C13 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C14 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C15 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C16 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C17 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.36fF
C18 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C19 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C20 7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C21 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C22 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C23 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.39fF
C24 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C25 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 m6_733_n10# 2.39fF
C26 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C27 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C28 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C29 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C30 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.36fF
C31 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C32 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C33 7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C34 D1 m6_733_n10# 38.89fF
C35 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C36 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C37 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C38 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C39 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 m6_733_n10# 2.39fF
C40 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C41 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C42 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C43 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C44 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.36fF
C45 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C46 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C47 7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C48 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C49 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C50 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.39fF
C51 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C52 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 m6_733_n10# 2.39fF
C53 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C54 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C55 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C56 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C57 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.36fF
C58 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C59 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C60 7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C61 7BitDac_0/6BitDac_1/V_out6 m6_733_n10# 2.06fF
C62 7BitDac_1/V_out7 m6_733_n10# 2.40fF
C63 VA m6_733_n10# 465.12fF
C64 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C65 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C66 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C67 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C68 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 m6_733_n10# 2.39fF
C69 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C70 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C71 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C72 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C73 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.36fF
C74 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C75 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C76 7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C77 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C78 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C79 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.39fF
C80 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C81 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 m6_733_n10# 2.39fF
C82 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C83 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C84 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C85 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C86 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.36fF
C87 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C88 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C89 7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C90 D0 m6_733_n10# 50.57fF
C91 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C92 D2 m6_733_n10# 30.50fF
C93 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C94 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C95 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C96 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 m6_733_n10# 2.39fF
C97 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C98 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C99 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C100 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C101 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.36fF
C102 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C103 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C104 7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C105 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C106 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C107 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.39fF
C108 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C109 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 m6_733_n10# 2.39fF
C110 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C111 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C112 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C113 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 m6_733_n10# 2.43fF
C114 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 m6_733_n10# 2.36fF
C115 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 m6_733_n10# 2.17fF
C116 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 m6_733_n10# 2.11fF
C117 7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 m6_733_n10# 2.35fF
C118 7BitDac_1/6BitDac_1/V_out6 m6_733_n10# 2.06fF



valpha  R_in8 Gnd 3.3
vbeta  VA Gnd 3.3
vzero D0 Gnd pulse(0 1.8 0.1m 60p 60p 0.1m 0.2m)
vone  D1 Gnd pulse(0 1.8 0.2m 60p 60p 0.2m 0.4m)
vtwo  D2 Gnd pulse(0 1.8 0.4m 60p 60p 0.4m 0.8m)
vthree D3 Gnd pulse(0 1.8 0.8m 60p 60p 0.8m 1.6m)
vfour D4 Gnd pulse (0 1.8 1.6m 60p 60p 1.6m 3.2m)
vfive D5 Gnd pulse (0 1.8 3.2m 60p 60p 3.2m 6.4m)
vsix D6 Gnd pulse (0 1.8 6.4m 60p 60p 6.4m 12.8m)
vseven D7 Gnd pulse (0 1.8 12.8m 60p 60p 12.8m 25.6m)

.tran 0.01m 25.6m
.control
run

plot V(V_out8) V(D0)

.endc
.end

