* SPICE3 file created from 5BitDac.ext - technology: scmos
.model polyResistor R ( TC1=0 TC2=0 RSH=7.7 DEFW=1.E-7 NARROW=0.0 TNOM=27)

.model pfet PMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=4.1589E17 VTH0=-0.3938813 K1=0.5479015 K2=0.0360586 K3=0.0993095 K3B=5.7086622 W0=1E-6 NLX=1.313191E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=0.4911363 DVT1=0.2227356 DVT2=0.1 U0=115.6852975 UA=1.505832E-9 UB=1E-21 UC=-1E-10 VSAT=1.329694E5 A0=1.7590478 AGS=0.3641621 B0=3.427126E-7 B1=1.062928E-6 KETA=0.0134667 A1=0.6859506 A2=0.3506788 RDSW=168.5705677 PRWG=0.5 PRWB=-0.4987371 WR=1 WINT=0 LINT=3.028832E-8 XL=0 XW=-1E-8 DWG=-2.349633E-8 DWB=-7.152486E-9 VOFF=-0.0994037 NFACTOR=1.9424315 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=0.0608072 ETAB=-0.0426148 DSUB=0.7343015 PCLM=3.2579974 PDIBLC1=7.229527E-6 PDIBLC2=0.025389 PDIBLCB=-1E-3 DROUT=0 PSCBE1=1.454878E10 PSCBE2=4.202027E-9 PVAG=15 DELTA=0.01 RSH=7.8 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=6.32E-10 CGSO=6.32E-10 CGBO=1E-12 CJ=1.172138E-3 PB=0.8421173 MJ=0.4109788 CJSW=2.242609E-10 PBSW=0.8 MJSW=0.3752089 CJSWG=4.22E-10 PBSWG=0.8 MJSWG=0.3752089 CF=0 PVTH0=1.888482E-3 PRDSW=11.5315407 PK2=1.559399E-3 WKETA=0.0319301 LKETA=2.955547E-3 PU0=-1.1105313 PUA=-4.62102E-11 PUB=1E-21 PVSAT=50 PETA0=1E-4 PKETA=-4.346368E-3)

.model nfet NMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=2.3549E17 VTH0=0.3823463 K1=0.5810697 K2=4.774618E-3 K3=0.0431669 K3B=1.1498346 W0=1E-7 NLX=1.910552E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=1.2894824 DVT1=0.3622063 DVT2=0.0713729 U0=280.633249 UA=-1.208537E-9 UB=2.158625E-18 UC=5.342807E-11 VSAT=9.366802E4 A0=1.7593146 AGS=0.3939741 B0=-6.413949E-9 B1=-1E-7 KETA=-5.180424E-4 A1=0 A2=1 RDSW=105.5517558 PRWG=0.5 PRWB=-0.1998871 WR=1 WINT=7.904732E-10 LINT=1.571424E-8 XL=0 XW=-1E-8 DWG=1.297221E-9 DWB=1.479041E-9 VOFF=-0.0955434 NFACTOR=2.4358891 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=3.104851E-3 ETAB=-2.512384E-5 DSUB=0.0167075 PCLM=0.8073191 PDIBLC1=0.1666161 PDIBLC2=3.112892E-3 PDIBLCB=-0.1 DROUT=0.7875618 PSCBE1=8E10 PSCBE2=9.213635E-10 PVAG=3.85243E-3 DELTA=0.01 RSH=6.7 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=7.08E-10 CGSO=7.08E-10 CGBO=1E-12 CJ=9.68858E-4 PB=0.8 MJ=0.3864502 CJSW=2.512138E-10 PBSW=0.809286 MJSW=0.1060414 CJSWG=3.3E-10 PBSWG=0.809286 MJSWG=0.1060414 CF=0 PVTH0=-1.192722E-3 PRDSW=-5 PK2=6.450505E-5 WKETA=-4.27294E-4 LKETA=-0.0104078 PU0=6.3268729 PUA=2.226552E-11 PUB=0 PVSAT=969.1480157 PETA0=1E-4 PKETA=-1.049509E-3)
.option scale=0.1u

M1000 switchNew_0/a_86_24# D4 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=4340 ps=2108
M1001 switchNew_0/a_105_20# switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1002 V_out5 switchNew_0/a_86_24# 4BitDac_0/V_out4 4BitDac_0/V_out4 pfet w=10 l=2
+  ad=140 pd=68 as=210 ps=102
M1003 4BitDac_0/V_out4 switchNew_0/a_105_20# V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=86 ps=64
M1004 switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=2205 ps=1512
M1005 switchNew_0/a_105_20# switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1006 V_out5 switchNew_0/a_86_24# 4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1007 V_out5 switchNew_0/a_105_20# 4BitDac_1/V_out4 V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1008 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1009 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1010 4BitDac_1/3BitDac_1/2BitDac_1/V_out2 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1011 4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1012 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1013 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1014 4BitDac_1/3BitDac_1/2BitDac_1/V_out2 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1015 4BitDac_1/3BitDac_1/2BitDac_1/V_out2 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1016 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1017 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1018 4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 4BitDac_1/3BitDac_1/2BitDac_1/gamma 4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1019 4BitDac_1/3BitDac_1/2BitDac_1/gamma 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1020 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1021 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1022 4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# gnd 4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=1558 ps=1522
R0 4BitDac_1/3BitDac_1/2BitDac_1/gamma gnd polyResistor w=2 l=62
R1 4BitDac_1/3BitDac_1/2BitDac_1/beta 4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
M1024 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1025 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1026 4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 4BitDac_1/3BitDac_1/2BitDac_1/alpha 4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1027 4BitDac_1/3BitDac_1/2BitDac_1/alpha 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1028 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1029 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1030 4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1031 4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_1/beta 4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R2 4BitDac_1/3BitDac_1/2BitDac_1/alpha 4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R3 4BitDac_1/3BitDac_1/2BitDac_0/delta 4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1032 4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1033 4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 4BitDac_1/3BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1034 4BitDac_1/3BitDac_1/V_out3 4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 4BitDac_1/3BitDac_1/2BitDac_0/V_out2 4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1035 4BitDac_1/3BitDac_1/2BitDac_0/V_out2 4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1036 4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1037 4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1038 4BitDac_1/3BitDac_1/V_out3 4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1039 4BitDac_1/3BitDac_1/V_out3 4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_1/V_out2 4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1041 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1042 4BitDac_1/3BitDac_1/2BitDac_0/V_out2 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1043 4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1044 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1045 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1046 4BitDac_1/3BitDac_1/2BitDac_0/V_out2 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1047 4BitDac_1/3BitDac_1/2BitDac_0/V_out2 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1048 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1049 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1050 4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 4BitDac_1/3BitDac_1/2BitDac_0/gamma 4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1051 4BitDac_1/3BitDac_1/2BitDac_0/gamma 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1052 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1053 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1054 4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1055 4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_0/delta 4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R4 4BitDac_1/3BitDac_1/2BitDac_0/gamma 4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
R5 4BitDac_1/3BitDac_1/2BitDac_0/beta 4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
M1056 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1057 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1058 4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 4BitDac_1/3BitDac_1/2BitDac_0/alpha 4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1059 4BitDac_1/3BitDac_1/2BitDac_0/alpha 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1060 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1061 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1062 4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1063 4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 4BitDac_1/3BitDac_1/2BitDac_0/beta 4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R6 4BitDac_1/3BitDac_1/2BitDac_0/alpha 4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R7 4BitDac_1/3BitDac_1/R_in3 4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1064 4BitDac_1/switchNew_0/a_86_24# D3 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1065 4BitDac_1/switchNew_0/a_105_20# 4BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1066 4BitDac_1/V_out4 4BitDac_1/switchNew_0/a_86_24# 4BitDac_1/3BitDac_0/V_out3 4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1067 4BitDac_1/3BitDac_0/V_out3 4BitDac_1/switchNew_0/a_105_20# 4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1068 4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1069 4BitDac_1/switchNew_0/a_105_20# 4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1070 4BitDac_1/V_out4 4BitDac_1/switchNew_0/a_86_24# 4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1071 4BitDac_1/V_out4 4BitDac_1/switchNew_0/a_105_20# 4BitDac_1/3BitDac_1/V_out3 4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1072 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1073 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1074 4BitDac_1/3BitDac_0/2BitDac_1/V_out2 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1075 4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1076 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1077 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1078 4BitDac_1/3BitDac_0/2BitDac_1/V_out2 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1079 4BitDac_1/3BitDac_0/2BitDac_1/V_out2 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1080 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1081 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1082 4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 4BitDac_1/3BitDac_0/2BitDac_1/gamma 4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1083 4BitDac_1/3BitDac_0/2BitDac_1/gamma 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1084 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1085 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1086 4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1087 4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 4BitDac_1/3BitDac_1/R_in3 4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R8 4BitDac_1/3BitDac_0/2BitDac_1/gamma 4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
R9 4BitDac_1/3BitDac_0/2BitDac_1/beta 4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
M1088 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1089 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1090 4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 4BitDac_1/3BitDac_0/2BitDac_1/alpha 4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1091 4BitDac_1/3BitDac_0/2BitDac_1/alpha 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1092 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1093 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1094 4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1095 4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_1/beta 4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R10 4BitDac_1/3BitDac_0/2BitDac_1/alpha 4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R11 4BitDac_1/3BitDac_0/2BitDac_0/delta 4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1096 4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1097 4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 4BitDac_1/3BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1098 4BitDac_1/3BitDac_0/V_out3 4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 4BitDac_1/3BitDac_0/2BitDac_0/V_out2 4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1099 4BitDac_1/3BitDac_0/2BitDac_0/V_out2 4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1100 4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1101 4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1102 4BitDac_1/3BitDac_0/V_out3 4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1103 4BitDac_1/3BitDac_0/V_out3 4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_1/V_out2 4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1104 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1105 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1106 4BitDac_1/3BitDac_0/2BitDac_0/V_out2 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1107 4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1108 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1109 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1110 4BitDac_1/3BitDac_0/2BitDac_0/V_out2 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1111 4BitDac_1/3BitDac_0/2BitDac_0/V_out2 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1112 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1113 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1114 4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 4BitDac_1/3BitDac_0/2BitDac_0/gamma 4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1115 4BitDac_1/3BitDac_0/2BitDac_0/gamma 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1116 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1117 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1118 4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1119 4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_0/delta 4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R12 4BitDac_1/3BitDac_0/2BitDac_0/gamma 4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
R13 4BitDac_1/3BitDac_0/2BitDac_0/beta 4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
M1120 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1121 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1122 4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 4BitDac_1/3BitDac_0/2BitDac_0/alpha 4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1123 4BitDac_1/3BitDac_0/2BitDac_0/alpha 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1124 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1125 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1126 4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1127 4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 4BitDac_1/3BitDac_0/2BitDac_0/beta 4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R14 4BitDac_1/3BitDac_0/2BitDac_0/alpha 4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R15 4BitDac_1/R_in4 4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1128 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1129 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1130 4BitDac_0/3BitDac_1/2BitDac_1/V_out2 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1131 4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1132 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1133 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1134 4BitDac_0/3BitDac_1/2BitDac_1/V_out2 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1135 4BitDac_0/3BitDac_1/2BitDac_1/V_out2 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1136 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1137 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1138 4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 4BitDac_0/3BitDac_1/2BitDac_1/gamma 4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1139 4BitDac_0/3BitDac_1/2BitDac_1/gamma 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1140 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1141 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1142 4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1143 4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 4BitDac_1/R_in4 4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R16 4BitDac_0/3BitDac_1/2BitDac_1/gamma 4BitDac_1/R_in4 polyResistor w=2 l=62
R17 4BitDac_0/3BitDac_1/2BitDac_1/beta 4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
M1144 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1145 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1146 4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 4BitDac_0/3BitDac_1/2BitDac_1/alpha 4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1147 4BitDac_0/3BitDac_1/2BitDac_1/alpha 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1148 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1149 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1150 4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1151 4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_1/beta 4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R18 4BitDac_0/3BitDac_1/2BitDac_1/alpha 4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R19 4BitDac_0/3BitDac_1/2BitDac_0/delta 4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1152 4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1153 4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 4BitDac_0/3BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1154 4BitDac_0/3BitDac_1/V_out3 4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 4BitDac_0/3BitDac_1/2BitDac_0/V_out2 4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1155 4BitDac_0/3BitDac_1/2BitDac_0/V_out2 4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1156 4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1157 4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1158 4BitDac_0/3BitDac_1/V_out3 4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 4BitDac_0/3BitDac_1/V_out3 4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_1/V_out2 4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1160 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1161 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1162 4BitDac_0/3BitDac_1/2BitDac_0/V_out2 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1163 4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1164 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1165 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1166 4BitDac_0/3BitDac_1/2BitDac_0/V_out2 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1167 4BitDac_0/3BitDac_1/2BitDac_0/V_out2 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1168 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1169 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1170 4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 4BitDac_0/3BitDac_1/2BitDac_0/gamma 4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1171 4BitDac_0/3BitDac_1/2BitDac_0/gamma 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1172 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1173 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1174 4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1175 4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_0/delta 4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R20 4BitDac_0/3BitDac_1/2BitDac_0/gamma 4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
R21 4BitDac_0/3BitDac_1/2BitDac_0/beta 4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
M1176 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1177 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1178 4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 4BitDac_0/3BitDac_1/2BitDac_0/alpha 4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1179 4BitDac_0/3BitDac_1/2BitDac_0/alpha 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1180 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1181 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1182 4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1183 4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 4BitDac_0/3BitDac_1/2BitDac_0/beta 4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R22 4BitDac_0/3BitDac_1/2BitDac_0/alpha 4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R23 4BitDac_0/3BitDac_1/R_in3 4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1184 4BitDac_0/switchNew_0/a_86_24# D3 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1185 4BitDac_0/switchNew_0/a_105_20# 4BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1186 4BitDac_0/V_out4 4BitDac_0/switchNew_0/a_86_24# 4BitDac_0/3BitDac_0/V_out3 4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1187 4BitDac_0/3BitDac_0/V_out3 4BitDac_0/switchNew_0/a_105_20# 4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1188 4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1189 4BitDac_0/switchNew_0/a_105_20# 4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1190 4BitDac_0/V_out4 4BitDac_0/switchNew_0/a_86_24# 4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1191 4BitDac_0/V_out4 4BitDac_0/switchNew_0/a_105_20# 4BitDac_0/3BitDac_1/V_out3 4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1193 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1194 4BitDac_0/3BitDac_0/2BitDac_1/V_out2 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1195 4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1196 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1197 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1198 4BitDac_0/3BitDac_0/2BitDac_1/V_out2 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1199 4BitDac_0/3BitDac_0/2BitDac_1/V_out2 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1200 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1201 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1202 4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 4BitDac_0/3BitDac_0/2BitDac_1/gamma 4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1203 4BitDac_0/3BitDac_0/2BitDac_1/gamma 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1204 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1205 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1206 4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1207 4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 4BitDac_0/3BitDac_1/R_in3 4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R24 4BitDac_0/3BitDac_0/2BitDac_1/gamma 4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
R25 4BitDac_0/3BitDac_0/2BitDac_1/beta 4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
M1208 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1209 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1210 4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 4BitDac_0/3BitDac_0/2BitDac_1/alpha 4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1211 4BitDac_0/3BitDac_0/2BitDac_1/alpha 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1212 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1213 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1214 4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1215 4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_1/beta 4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R26 4BitDac_0/3BitDac_0/2BitDac_1/alpha 4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R27 4BitDac_0/3BitDac_0/2BitDac_0/delta 4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1216 4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1217 4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 4BitDac_0/3BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1218 4BitDac_0/3BitDac_0/V_out3 4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 4BitDac_0/3BitDac_0/2BitDac_0/V_out2 4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1219 4BitDac_0/3BitDac_0/2BitDac_0/V_out2 4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1220 4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1221 4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1222 4BitDac_0/3BitDac_0/V_out3 4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 4BitDac_0/3BitDac_0/V_out3 4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_1/V_out2 4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1224 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1225 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1226 4BitDac_0/3BitDac_0/2BitDac_0/V_out2 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1227 4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1228 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1229 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1230 4BitDac_0/3BitDac_0/2BitDac_0/V_out2 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1231 4BitDac_0/3BitDac_0/2BitDac_0/V_out2 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1232 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1233 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1234 4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 4BitDac_0/3BitDac_0/2BitDac_0/gamma 4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1235 4BitDac_0/3BitDac_0/2BitDac_0/gamma 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1236 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1237 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1238 4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1239 4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_0/delta 4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R28 4BitDac_0/3BitDac_0/2BitDac_0/gamma 4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
R29 4BitDac_0/3BitDac_0/2BitDac_0/beta 4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
M1240 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1241 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1242 4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 4BitDac_0/3BitDac_0/2BitDac_0/alpha 4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1243 4BitDac_0/3BitDac_0/2BitDac_0/alpha 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1244 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1245 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1246 4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1247 4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 4BitDac_0/3BitDac_0/2BitDac_0/beta 4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R30 4BitDac_0/3BitDac_0/2BitDac_0/alpha 4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R31 R_in5 4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
C0 D2 D1 5.43fF
C1 4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.17fF
C2 4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C3 4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C4 4BitDac_0/3BitDac_1/V_out3 gnd 2.22fF
C5 4BitDac_0/V_out4 gnd 2.30fF
C6 4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.17fF
C7 4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C8 D1 gnd 2.85fF
C9 4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.17fF
C10 4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C11 4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C12 4BitDac_1/3BitDac_1/V_out3 gnd 2.22fF
C13 D0 gnd 5.07fF
C14 4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.17fF
C15 4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C16 Vdd gnd 29.90fF





valpha  R_in5 Gnd 3.3
vbeta  Vdd Gnd 3.3
vzero D0 Gnd pulse(0 1.8 0.1m 60p 60p 0.1m 0.2m)
vone  D1 Gnd pulse(0 1.8 0.2m 60p 60p 0.2m 0.4m)
vtwo  D2 Gnd pulse(0 1.8 0.4m 60p 60p 0.4m 0.8m)
vthree D3 Gnd pulse(0 1.8 0.8m 60p 60p 0.8m 1.6m)
vfour D4 Gnd pulse (0 1.8 1.6m 60p 60p 1.6m 3.2m)
.tran 0.01m 3.2m
.control
run

plot V(V_out5) V(D0)

.endc
.end







