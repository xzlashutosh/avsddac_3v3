* E:\esim-DAC\2_bit_dac\2_bit_dac.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 08/12/20 07:10:50

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  Net-_R1-Pad2_ GND 3.3		
R1  Net-_R1-Pad1_ Net-_R1-Pad2_ 250		
R2  Net-_R2-Pad1_ Net-_R1-Pad1_ 250		
R3  Net-_R3-Pad1_ Net-_R2-Pad1_ 250		
R4  GND Net-_R3-Pad1_ 250		
v3  Vtwo GND pulse		
v2  Vone GND pulse		
U1  Voutput plot_v1		
U2  Vone plot_v2		
X1  Vone Net-_R1-Pad1_ Net-_R2-Pad1_ /vmid1 switch		
X2  Vone Net-_R3-Pad1_ GND /vmid2 switch		
X3  Vtwo /vmid1 /vmid2 Voutput switch		
C1  Voutput GND 5p		

.end
