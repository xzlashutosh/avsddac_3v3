* C:\FOSSEE\eSim\library\SubcircuitLibrary\3_bit_dac\3_bit_dac.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 08/12/20 14:07:00

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad3_ Net-_X1-Pad2_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_X1-Pad5_ 2_bit_dac		
X2  Net-_X1-Pad2_ Net-_U1-Pad4_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_X2-Pad5_ 2_bit_dac		
X3  Net-_U1-Pad5_ Net-_X1-Pad5_ Net-_X2-Pad5_ Net-_U1-Pad6_ switch		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ PORT		

.end
