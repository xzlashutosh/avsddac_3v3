magic
tech scmos
timestamp 1599268620
<< metal1 >>
rect -7 210 -2 216
rect 272 95 286 98
rect 283 49 286 95
rect 212 45 286 49
rect 212 37 215 45
rect -9 14 13 20
rect 157 1 162 5
rect 272 4 283 7
rect 209 -38 212 -22
rect 209 -42 290 -38
rect 287 -94 290 -42
rect 270 -97 290 -94
rect 7 -182 11 -178
<< metal3 >>
rect 17 202 21 210
rect 152 150 156 159
rect 136 92 154 97
rect 16 49 20 56
rect 16 5 19 49
rect 136 -30 140 92
rect 136 -34 154 -30
rect 150 -43 154 -34
<< metal5 >>
rect 80 94 101 99
rect 96 88 133 94
rect 96 1 101 88
rect 128 62 133 88
rect 128 59 170 62
rect 166 49 170 59
rect 166 48 180 49
rect 166 45 188 48
rect 176 44 188 45
<< metal6 >>
rect 24 -87 33 14
rect 175 -37 181 -32
rect 160 -44 181 -37
rect 160 -140 165 -44
use 2BitDac  2BitDac_0
timestamp 1599268620
transform 1 0 -61 0 1 183
box 52 -171 333 27
use switchNew  switchNew_0
timestamp 1599222484
transform 1 0 85 0 1 -35
box 69 -1 187 81
use 2BitDac  2BitDac_1
timestamp 1599268620
transform 1 0 -63 0 1 -9
box 52 -171 333 27
<< labels >>
rlabel metal1 283 4 283 7 7 V_out3
rlabel metal1 -7 216 -2 216 5 R_in3
rlabel metal1 7 -182 11 -182 1 R_out3
<< end >>
