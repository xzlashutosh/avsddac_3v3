magic
tech scmos
timestamp 1599268620
<< metal1 >>
rect -2 403 3 404
rect 287 191 301 194
rect 298 42 301 191
rect 213 39 301 42
rect 213 20 216 39
rect -6 0 16 5
rect 162 -17 163 -13
rect 273 -14 299 -11
rect 209 -53 213 -44
rect 209 -56 293 -53
rect 290 -205 293 -56
rect 283 -208 293 -205
rect 8 -395 12 -394
<< m2contact >>
rect 162 187 166 195
rect 156 -212 165 -204
<< m3contact >>
rect 162 187 166 195
rect 156 -212 165 -204
<< metal3 >>
rect 22 397 26 401
rect 157 346 161 358
rect 167 245 170 339
rect 162 242 170 245
rect 162 195 165 242
rect 162 100 165 187
rect 162 95 173 100
rect 144 91 158 92
rect 138 87 158 91
rect 159 87 160 91
rect 20 3 24 49
rect 18 0 24 3
rect 18 -9 22 0
rect 138 -57 142 87
rect 168 84 173 95
rect 162 79 173 84
rect 138 -60 157 -57
rect 162 -109 165 79
rect 162 -112 166 -109
rect 163 -113 166 -112
rect 163 -124 167 -113
rect 162 -127 167 -124
rect 162 -204 165 -127
<< metal5 >>
rect 118 95 125 96
rect 79 89 125 95
rect 118 28 125 89
rect 118 23 189 28
rect 118 -18 125 23
<< metal6 >>
rect 72 -104 77 12
rect 177 -60 182 -48
rect 177 -65 206 -60
rect 51 -109 77 -104
rect 201 -155 206 -65
rect 173 -160 206 -155
use 3BitDac  3BitDac_0
timestamp 1599268620
transform 1 0 5 0 1 187
box -11 -182 290 216
use switchNew  switchNew_0
timestamp 1599222484
transform 1 0 86 0 1 -53
box 69 -1 187 81
use 3BitDac  3BitDac_1
timestamp 1599268620
transform 1 0 1 0 1 -212
box -11 -182 290 216
<< labels >>
rlabel metal1 299 -14 299 -11 7 V_out4
rlabel metal1 -2 404 3 404 5 R_in4
rlabel metal1 8 -395 12 -395 1 R_out4
<< end >>
