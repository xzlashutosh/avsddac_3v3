* D:\DAC\esim-DAC\10_bit_dac\10_bit_dac.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 08/22/20 13:05:10

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v9  Net-_X1-Pad9_ GND 3.3		
X3  Net-_X3-Pad1_ Net-_X1-Pad12_ Net-_X2-Pad12_ Vout switch		
v1  Net-_X1-Pad1_ GND pulse		
v2  Net-_X1-Pad2_ GND pulse		
v3  Net-_X1-Pad3_ GND pulse		
v4  Net-_X1-Pad4_ GND pulse		
v5  Net-_X1-Pad5_ GND pulse		
v11  Net-_X3-Pad1_ GND pulse		
U1  Vout plot_v1		
v6  Net-_X1-Pad6_ GND pulse		
v7  Net-_X1-Pad7_ GND pulse		
v8  Net-_X1-Pad8_ GND pulse		
v10  Net-_X1-Pad11_ GND pulse		
X1  Net-_X1-Pad1_ Net-_X1-Pad2_ Net-_X1-Pad3_ Net-_X1-Pad4_ Net-_X1-Pad5_ Net-_X1-Pad6_ Net-_X1-Pad7_ Net-_X1-Pad8_ Net-_X1-Pad9_ Net-_X1-Pad10_ Net-_X1-Pad11_ Net-_X1-Pad12_ 9_bit_dac		
X2  Net-_X1-Pad1_ Net-_X1-Pad2_ Net-_X1-Pad3_ Net-_X1-Pad4_ Net-_X1-Pad5_ Net-_X1-Pad6_ Net-_X1-Pad7_ Net-_X1-Pad8_ Net-_X1-Pad10_ GND Net-_X1-Pad11_ Net-_X2-Pad12_ 9_bit_dac		
C1  Vout GND 5000p		

.end
