* SPICE3 file created from 9BitDac.ext - technology: scmos


.model polyResistor R ( TC1=0 TC2=0 RSH=7.7 DEFW=1.E-7 NARROW=0.0 TNOM=27)

.model pfet PMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=4.1589E17 VTH0=-0.3938813 K1=0.5479015 K2=0.0360586 K3=0.0993095 K3B=5.7086622 W0=1E-6 NLX=1.313191E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=0.4911363 DVT1=0.2227356 DVT2=0.1 U0=115.6852975 UA=1.505832E-9 UB=1E-21 UC=-1E-10 VSAT=1.329694E5 A0=1.7590478 AGS=0.3641621 B0=3.427126E-7 B1=1.062928E-6 KETA=0.0134667 A1=0.6859506 A2=0.3506788 RDSW=168.5705677 PRWG=0.5 PRWB=-0.4987371 WR=1 WINT=0 LINT=3.028832E-8 XL=0 XW=-1E-8 DWG=-2.349633E-8 DWB=-7.152486E-9 VOFF=-0.0994037 NFACTOR=1.9424315 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=0.0608072 ETAB=-0.0426148 DSUB=0.7343015 PCLM=3.2579974 PDIBLC1=7.229527E-6 PDIBLC2=0.025389 PDIBLCB=-1E-3 DROUT=0 PSCBE1=1.454878E10 PSCBE2=4.202027E-9 PVAG=15 DELTA=0.01 RSH=7.8 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=6.32E-10 CGSO=6.32E-10 CGBO=1E-12 CJ=1.172138E-3 PB=0.8421173 MJ=0.4109788 CJSW=2.242609E-10 PBSW=0.8 MJSW=0.3752089 CJSWG=4.22E-10 PBSWG=0.8 MJSWG=0.3752089 CF=0 PVTH0=1.888482E-3 PRDSW=11.5315407 PK2=1.559399E-3 WKETA=0.0319301 LKETA=2.955547E-3 PU0=-1.1105313 PUA=-4.62102E-11 PUB=1E-21 PVSAT=50 PETA0=1E-4 PKETA=-4.346368E-3)

.model nfet NMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=2.3549E17 VTH0=0.3823463 K1=0.5810697 K2=4.774618E-3 K3=0.0431669 K3B=1.1498346 W0=1E-7 NLX=1.910552E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=1.2894824 DVT1=0.3622063 DVT2=0.0713729 U0=280.633249 UA=-1.208537E-9 UB=2.158625E-18 UC=5.342807E-11 VSAT=9.366802E4 A0=1.7593146 AGS=0.3939741 B0=-6.413949E-9 B1=-1E-7 KETA=-5.180424E-4 A1=0 A2=1 RDSW=105.5517558 PRWG=0.5 PRWB=-0.1998871 WR=1 WINT=7.904732E-10 LINT=1.571424E-8 XL=0 XW=-1E-8 DWG=1.297221E-9 DWB=1.479041E-9 VOFF=-0.0955434 NFACTOR=2.4358891 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=3.104851E-3 ETAB=-2.512384E-5 DSUB=0.0167075 PCLM=0.8073191 PDIBLC1=0.1666161 PDIBLC2=3.112892E-3 PDIBLCB=-0.1 DROUT=0.7875618 PSCBE1=8E10 PSCBE2=9.213635E-10 PVAG=3.85243E-3 DELTA=0.01 RSH=6.7 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=7.08E-10 CGSO=7.08E-10 CGBO=1E-12 CJ=9.68858E-4 PB=0.8 MJ=0.3864502 CJSW=2.512138E-10 PBSW=0.809286 MJSW=0.1060414 CJSWG=3.3E-10 PBSWG=0.809286 MJSWG=0.1060414 CF=0 PVTH0=-1.192722E-3 PRDSW=-5 PK2=6.450505E-5 WKETA=-4.27294E-4 LKETA=-0.0104078 PU0=6.3268729 PUA=2.226552E-11 PUB=0 PVSAT=969.1480157 PETA0=1E-4 PKETA=-1.049509E-3)



.option scale=0.1u

M1000 8BitDac_1/7BitDac_1/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=71540 ps=34748
M1001 8BitDac_1/7BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1002 8BitDac_1/7BitDac_1/V_out7 8BitDac_1/7BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/V_out6 8BitDac_1/7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1003 8BitDac_1/7BitDac_1/6BitDac_0/V_out6 8BitDac_1/7BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/V_out7 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1004 8BitDac_1/7BitDac_1/switchNew_0/a_86_24# D6 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=35805 ps=24552
M1005 8BitDac_1/7BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1006 8BitDac_1/7BitDac_1/V_out7 8BitDac_1/7BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1007 8BitDac_1/7BitDac_1/V_out7 8BitDac_1/7BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/V_out6 8BitDac_1/7BitDac_1/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1008 8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1009 8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1010 8BitDac_1/7BitDac_1/6BitDac_1/V_out6 8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1011 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1012 8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1013 8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1014 8BitDac_1/7BitDac_1/6BitDac_1/V_out6 8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1015 8BitDac_1/7BitDac_1/6BitDac_1/V_out6 8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 8BitDac_1/7BitDac_1/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1016 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1017 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1018 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1019 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1020 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1021 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1022 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1023 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1024 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1025 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1026 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1027 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1028 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1029 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1030 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1031 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1032 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1033 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1034 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1035 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1036 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1037 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1038 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1039 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# gnd 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=24598 ps=24562
R0 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma gnd polyResistor w=2 l=62
M1040 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1041 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1042 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1043 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1044 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1045 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1046 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1047 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1048 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1049 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1050 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1051 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1052 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1053 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1054 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1057 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1058 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1059 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1060 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1061 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1062 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1063 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1064 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1065 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1066 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1067 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1068 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1069 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1070 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1071 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1072 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1073 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1074 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1075 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1076 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1077 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1078 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1079 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R5 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R6 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R7 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1080 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1081 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1082 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1083 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1084 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1085 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1086 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1089 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1090 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1091 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1092 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1093 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1094 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1095 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1096 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1097 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1098 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1099 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1100 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1101 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1102 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1103 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R8 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M1104 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1105 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1106 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1107 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1108 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1109 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1110 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1111 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R9 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R10 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R11 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1112 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1113 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1114 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1115 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1116 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1117 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1118 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1121 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1122 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1123 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1124 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1125 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1126 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1127 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1128 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1129 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1130 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1131 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1132 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1133 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1134 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1135 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R12 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1136 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1137 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1138 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1139 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1140 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1141 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1142 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1143 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R13 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R14 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R15 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1144 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1145 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1146 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1147 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1148 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1149 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1150 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1151 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1152 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1153 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1154 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1155 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1156 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1157 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1158 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1159 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R16 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M1160 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1161 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1162 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1163 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1164 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1165 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1166 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1167 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R17 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R18 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R19 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1168 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1169 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1170 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1171 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1172 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1173 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1174 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1177 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1178 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1179 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1180 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1181 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1182 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1183 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1184 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1185 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1186 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1187 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1188 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1189 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1190 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1191 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R20 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1192 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1193 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1194 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1195 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1196 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1197 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1198 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1199 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R21 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R22 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R23 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1200 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1201 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1202 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1203 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1204 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1205 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1206 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1209 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1210 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1211 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1212 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1213 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1214 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1215 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1216 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1217 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1218 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1219 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1220 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1221 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1222 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1223 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R24 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M1224 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1225 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1226 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1227 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1228 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1229 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1230 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1231 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R25 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R26 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R27 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1232 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1233 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1234 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1235 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1236 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1237 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1238 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1240 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1241 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1242 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1243 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1244 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1245 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1246 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1247 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1248 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1249 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1250 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1251 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1252 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1253 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1254 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1255 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R28 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1256 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1257 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1258 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1259 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1260 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1261 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1262 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1263 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R29 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R30 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R31 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1264 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1265 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1266 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1267 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1268 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1269 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1270 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1271 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1272 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1273 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1274 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1275 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1276 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1277 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1278 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1279 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1280 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1281 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1282 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1283 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1284 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1285 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1286 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1287 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R32 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M1288 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1289 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1290 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1291 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1292 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1293 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1294 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1295 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R33 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R34 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R35 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1296 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1297 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1298 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1299 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1300 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1301 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1302 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1303 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1304 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1305 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1306 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1307 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1308 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1309 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1310 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1311 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1312 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1313 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1314 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1315 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1316 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1317 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1318 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1319 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R36 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1320 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1321 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1322 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1323 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1324 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1325 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1326 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1327 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R37 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R38 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R39 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1328 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1329 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1330 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1331 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1332 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1333 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1334 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1335 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1336 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1337 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1338 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1339 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1340 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1341 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1342 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1343 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1344 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1345 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1346 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1347 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1348 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1349 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1350 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1351 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R40 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M1352 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1353 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1354 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1355 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1356 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1357 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1358 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1359 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R41 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R42 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R43 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1360 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1361 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1362 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1363 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1364 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1365 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1366 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1367 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1368 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1369 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1370 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1371 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1372 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1373 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1374 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1375 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1376 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1377 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1378 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1379 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1380 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1381 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1382 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1383 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R44 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1384 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1385 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1386 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1387 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1388 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1389 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1390 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1391 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R45 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R46 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R47 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1392 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1393 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1394 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1395 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1396 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1397 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1398 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1399 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1400 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1401 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1402 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1403 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1404 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1405 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1406 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1407 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R48 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M1408 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1409 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1410 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1411 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1412 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1413 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1414 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1415 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R49 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R50 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R51 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1416 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1417 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1418 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1419 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1420 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1421 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1422 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1423 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1424 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1425 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1426 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1427 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1428 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1429 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1430 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1431 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1432 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1433 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1434 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1435 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1436 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1437 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1438 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1439 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R52 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1440 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1441 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1442 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1443 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1444 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1445 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1446 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1447 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R53 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R54 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R55 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1448 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1449 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1450 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1451 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1452 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1453 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1454 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1455 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1456 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1457 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1458 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1459 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1460 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1461 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1462 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1463 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1464 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1465 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1466 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1467 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1468 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1469 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1470 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1471 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R56 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M1472 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1473 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1474 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1475 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1476 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1477 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1478 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1479 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R57 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R58 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R59 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1480 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1481 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1482 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1483 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1484 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1485 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1486 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1487 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1488 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1489 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1490 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1491 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1492 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1493 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1494 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1495 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1496 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1497 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1498 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1499 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1500 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1501 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1502 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1503 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R60 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1504 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1505 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1506 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1507 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1508 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1509 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1510 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1511 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R61 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R62 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R63 8BitDac_1/7BitDac_1/6BitDac_1/R_in6 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1512 8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1513 8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1514 8BitDac_1/7BitDac_1/6BitDac_0/V_out6 8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1515 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1516 8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1517 8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1518 8BitDac_1/7BitDac_1/6BitDac_0/V_out6 8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1519 8BitDac_1/7BitDac_1/6BitDac_0/V_out6 8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 8BitDac_1/7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1520 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1521 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1522 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1523 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1524 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1525 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1526 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1527 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1528 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1529 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1530 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1531 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1532 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1533 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1534 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1535 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1536 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1537 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1538 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1539 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1540 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1541 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1542 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_1/R_in6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1543 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_1/R_in6 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R64 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_1/R_in6 polyResistor w=2 l=62
M1544 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1545 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1546 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1547 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1548 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1549 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1550 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1551 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R65 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R66 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R67 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1552 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1553 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1554 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1555 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1556 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1557 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1558 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1559 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1560 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1561 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1562 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1563 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1564 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1565 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1566 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1567 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1568 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1569 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1570 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1571 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1572 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1573 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1574 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1575 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R68 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1576 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1577 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1578 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1579 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1580 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1581 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1582 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1583 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R69 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R70 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R71 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1584 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1585 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1586 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1587 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1588 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1589 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1590 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1591 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1592 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1593 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1594 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1595 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1596 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1597 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1598 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1599 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1600 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1601 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1602 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1603 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1604 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1605 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1606 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1607 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R72 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M1608 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1609 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1610 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1611 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1612 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1613 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1614 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1615 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R73 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R74 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R75 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1616 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1617 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1618 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1619 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1620 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1621 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1622 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1623 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1624 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1625 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1626 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1627 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1628 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1629 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1630 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1631 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1632 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1633 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1634 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1635 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1636 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1637 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1638 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1639 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R76 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1640 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1641 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1642 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1643 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1644 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1645 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1646 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1647 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R77 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R78 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R79 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1648 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1649 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1650 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1651 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1652 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1653 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1654 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1655 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1656 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1657 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1658 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1659 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1660 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1661 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1662 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1663 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R80 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M1664 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1665 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1666 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1667 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1668 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1669 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1670 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1671 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R81 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R82 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R83 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1672 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1673 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1674 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1675 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1676 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1677 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1678 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1679 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1680 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1681 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1682 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1683 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1684 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1685 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1686 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1687 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1688 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1689 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1690 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1691 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1692 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1693 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1694 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1695 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R84 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1696 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1697 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1698 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1699 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1700 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1701 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1702 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1703 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R85 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R86 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R87 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1704 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1705 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1706 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1707 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1708 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1709 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1710 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1711 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1712 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1713 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1714 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1715 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1716 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1717 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1718 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1719 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1720 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1721 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1722 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1723 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1724 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1725 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1726 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1727 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R88 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M1728 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1729 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1730 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1731 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1732 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1733 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1734 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1735 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R89 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R90 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R91 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1736 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1737 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1738 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1739 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1740 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1741 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1742 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1743 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1744 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1745 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1746 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1747 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1748 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1749 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1750 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1751 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1752 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1753 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1754 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1755 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1756 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1757 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1758 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1759 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R92 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1760 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1761 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1762 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1763 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1764 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1765 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1766 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1767 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R93 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R94 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R95 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1768 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1769 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1770 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1771 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1772 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1773 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1774 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1775 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1776 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1777 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1778 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1779 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1780 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1781 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1782 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1783 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1784 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1785 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1786 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1787 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1788 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1789 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1790 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1791 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R96 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M1792 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1793 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1794 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1795 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1796 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1797 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1798 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1799 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R97 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R98 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R99 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1800 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1801 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1802 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1803 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1804 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1805 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1806 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1807 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1808 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1809 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1810 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1811 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1812 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1813 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1814 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1815 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1816 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1817 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1818 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1819 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1820 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1821 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1822 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1823 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R100 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1824 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1825 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1826 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1827 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1828 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1829 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1830 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1831 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R101 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R102 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R103 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1832 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1833 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1834 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1835 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1836 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1837 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1838 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1839 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1840 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1841 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1842 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1843 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1844 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1845 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1846 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1847 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1848 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1849 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1850 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1851 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1852 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1853 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1854 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1855 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R104 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M1856 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1857 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1858 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1859 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1860 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1861 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1862 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1863 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R105 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R106 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R107 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1864 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1865 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1866 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1867 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1868 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1869 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1870 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1871 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1872 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1873 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1874 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1875 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1876 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1877 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1878 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1879 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1880 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1881 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1882 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1883 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1884 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1885 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1886 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1887 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R108 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1888 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1889 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1890 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1891 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1892 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1893 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1894 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1895 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R109 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R110 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R111 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1896 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1897 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1898 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1899 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1900 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1901 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1902 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1903 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1904 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1905 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1906 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1907 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1908 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1909 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1910 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1911 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R112 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M1912 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1913 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1914 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1915 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1916 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1917 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1918 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1919 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R113 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R114 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R115 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1920 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1921 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1922 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1923 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1924 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1925 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1926 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1927 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1928 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1929 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1930 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1931 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1932 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1933 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1934 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1935 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1936 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1937 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1938 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1939 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1940 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1941 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1942 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1943 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R116 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1944 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1945 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1946 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1947 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1948 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1949 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1950 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1951 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R117 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R118 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R119 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1952 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1953 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1954 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1955 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1956 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1957 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1958 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1959 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1960 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1961 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1962 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1963 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1964 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1965 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1966 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1967 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1968 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1969 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1970 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1971 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1972 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1973 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1974 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1975 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R120 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M1976 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1977 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1978 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1979 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1980 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1981 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1982 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1983 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R121 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R122 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R123 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1984 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1985 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1986 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1987 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1988 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1989 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1990 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1991 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1992 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1993 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1994 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1995 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1996 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1997 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1998 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1999 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2000 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2001 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2002 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2003 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2004 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2005 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2006 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2007 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R124 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2008 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2009 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2010 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2011 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2012 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2013 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2014 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2015 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R125 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R126 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R127 8BitDac_1/7BitDac_1/R_in7 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2016 8BitDac_1/switchNew_0/a_86_24# D7 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2017 8BitDac_1/switchNew_0/a_105_21# 8BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2018 8BitDac_1/V_out8 8BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/V_out7 8BitDac_1/7BitDac_0/V_out7 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2019 8BitDac_1/7BitDac_0/V_out7 8BitDac_1/switchNew_0/a_105_21# 8BitDac_1/V_out8 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2020 8BitDac_1/switchNew_0/a_86_24# D7 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2021 8BitDac_1/switchNew_0/a_105_21# 8BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2022 8BitDac_1/V_out8 8BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_1/V_out7 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2023 8BitDac_1/V_out8 8BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_1/V_out7 8BitDac_1/V_out8 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2024 8BitDac_1/7BitDac_0/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2025 8BitDac_1/7BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2026 8BitDac_1/7BitDac_0/V_out7 8BitDac_1/7BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/V_out6 8BitDac_1/7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2027 8BitDac_1/7BitDac_0/6BitDac_0/V_out6 8BitDac_1/7BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/V_out7 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2028 8BitDac_1/7BitDac_0/switchNew_0/a_86_24# D6 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2029 8BitDac_1/7BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2030 8BitDac_1/7BitDac_0/V_out7 8BitDac_1/7BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2031 8BitDac_1/7BitDac_0/V_out7 8BitDac_1/7BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/V_out6 8BitDac_1/7BitDac_0/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2032 8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2033 8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2034 8BitDac_1/7BitDac_0/6BitDac_1/V_out6 8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2035 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2036 8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2037 8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2038 8BitDac_1/7BitDac_0/6BitDac_1/V_out6 8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2039 8BitDac_1/7BitDac_0/6BitDac_1/V_out6 8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 8BitDac_1/7BitDac_0/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2040 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2041 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2042 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2043 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2044 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2045 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2046 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2047 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2048 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2049 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2050 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2051 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2052 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2053 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2054 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2055 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2056 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2057 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2058 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2059 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2060 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2061 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2062 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_1/R_in7 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2063 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_1/R_in7 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R128 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_1/R_in7 polyResistor w=2 l=62
M2064 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2065 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2066 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2067 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2068 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2069 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2070 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2071 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R129 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R130 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R131 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2072 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2073 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2074 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2075 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2076 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2077 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2078 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2079 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2080 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2081 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2082 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2083 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2084 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2085 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2086 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2087 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2088 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2089 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2090 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2091 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2092 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2093 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2094 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2095 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R132 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2096 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2097 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2098 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2099 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2100 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2101 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2102 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2103 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R133 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R134 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R135 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2104 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2105 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2106 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2107 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2108 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2109 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2110 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2111 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2112 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2113 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2114 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2115 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2116 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2117 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2118 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2119 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2120 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2121 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2122 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2123 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2124 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2125 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2126 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2127 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R136 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M2128 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2129 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2130 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2131 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2132 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2133 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2134 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2135 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R137 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R138 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R139 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2136 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2137 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2138 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2139 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2140 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2141 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2142 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2143 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2144 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2145 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2146 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2147 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2148 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2149 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2150 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2151 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2152 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2153 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2154 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2155 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2156 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2157 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2158 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2159 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R140 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2160 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2161 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2162 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2163 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2164 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2165 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2166 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2167 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R141 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R142 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R143 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2168 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2169 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2170 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2171 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2172 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2173 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2174 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2175 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2176 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2177 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2178 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2179 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2180 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2181 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2182 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2183 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R144 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M2184 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2185 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2186 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2187 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2188 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2189 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2190 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2191 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R145 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R146 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R147 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2192 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2193 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2194 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2195 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2196 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2197 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2198 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2199 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2200 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2201 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2202 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2203 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2204 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2205 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2206 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2207 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2208 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2209 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2210 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2211 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2212 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2213 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2214 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2215 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R148 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2216 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2217 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2218 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2219 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2220 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2221 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2222 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2223 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R149 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R150 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R151 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2224 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2225 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2226 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2227 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2228 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2229 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2230 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2231 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2232 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2233 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2234 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2235 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2236 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2237 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2238 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2239 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2240 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2241 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2242 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2243 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2244 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2245 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2246 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2247 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R152 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M2248 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2249 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2250 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2251 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2252 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2253 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2254 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2255 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R153 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R154 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R155 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2256 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2257 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2258 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2259 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2260 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2261 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2262 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2263 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2264 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2265 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2266 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2267 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2268 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2269 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2270 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2271 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2272 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2273 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2274 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2275 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2276 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2277 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2278 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2279 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R156 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2280 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2281 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2282 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2283 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2284 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2285 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2286 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2287 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R157 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R158 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R159 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2288 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2289 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2290 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2291 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2292 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2293 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2294 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2295 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2296 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2297 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2298 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2299 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2300 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2301 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2302 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2303 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2304 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2305 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2306 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2307 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2308 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2309 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2310 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2311 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R160 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M2312 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2313 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2314 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2315 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2316 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2317 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2318 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2319 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R161 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R162 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R163 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2320 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2321 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2322 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2323 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2324 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2325 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2326 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2327 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2328 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2329 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2330 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2331 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2332 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2333 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2334 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2335 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2336 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2337 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2338 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2339 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2340 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2341 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2342 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2343 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R164 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2344 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2345 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2346 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2347 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2348 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2349 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2350 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2351 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R165 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R166 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R167 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2352 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2353 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2354 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2355 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2356 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2357 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2358 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2359 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2360 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2361 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2362 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2363 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2364 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2365 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2366 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2367 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2368 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2369 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2370 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2371 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2372 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2373 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2374 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2375 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R168 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M2376 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2377 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2378 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2379 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2380 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2381 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2382 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2383 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R169 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R170 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R171 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2384 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2385 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2386 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2387 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2388 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2389 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2390 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2391 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2392 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2393 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2394 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2395 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2396 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2397 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2398 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2399 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2400 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2401 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2402 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2403 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2404 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2405 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2406 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2407 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R172 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2408 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2409 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2410 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2411 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2412 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2413 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2414 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2415 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R173 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R174 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R175 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2416 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2417 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2418 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2419 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2420 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2421 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2422 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2423 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2424 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2425 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2426 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2427 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2428 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2429 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2430 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2431 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R176 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M2432 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2433 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2434 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2435 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2436 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2437 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2438 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2439 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R177 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R178 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R179 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2440 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2441 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2442 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2443 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2444 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2445 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2446 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2447 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2448 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2449 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2450 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2451 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2452 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2453 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2454 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2455 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2456 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2457 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2458 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2459 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2460 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2461 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2462 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2463 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R180 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2464 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2465 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2466 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2467 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2468 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2469 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2470 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2471 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R181 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R182 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R183 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2472 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2473 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2474 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2475 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2476 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2477 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2478 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2479 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2480 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2481 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2482 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2483 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2484 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2485 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2486 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2487 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2488 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2489 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2490 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2491 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2492 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2493 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2494 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2495 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R184 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M2496 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2497 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2498 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2499 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2500 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2501 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2502 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2503 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R185 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R186 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R187 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2504 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2505 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2506 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2507 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2508 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2509 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2510 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2511 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2512 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2513 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2514 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2515 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2516 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2517 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2518 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2519 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2520 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2521 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2522 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2523 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2524 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2525 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2526 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2527 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R188 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2528 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2529 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2530 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2531 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2532 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2533 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2534 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2535 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R189 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R190 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R191 8BitDac_1/7BitDac_0/6BitDac_1/R_in6 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2536 8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2537 8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2538 8BitDac_1/7BitDac_0/6BitDac_0/V_out6 8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2539 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2540 8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2541 8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2542 8BitDac_1/7BitDac_0/6BitDac_0/V_out6 8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2543 8BitDac_1/7BitDac_0/6BitDac_0/V_out6 8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 8BitDac_1/7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2544 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2545 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2546 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2547 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2548 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2549 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2550 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2551 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2552 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2553 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2554 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2555 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2556 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2557 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2558 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2559 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2560 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2561 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2562 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2563 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2564 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2565 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2566 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_1/R_in6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2567 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_1/R_in6 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R192 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_1/R_in6 polyResistor w=2 l=62
M2568 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2569 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2570 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2571 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2572 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2573 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2574 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2575 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R193 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R194 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R195 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2576 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2577 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2578 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2579 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2580 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2581 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2582 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2583 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2584 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2585 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2586 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2587 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2588 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2589 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2590 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2591 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2592 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2593 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2594 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2595 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2596 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2597 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2598 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2599 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R196 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2600 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2601 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2602 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2603 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2604 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2605 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2606 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2607 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R197 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R198 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R199 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2608 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2609 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2610 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2611 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2612 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2613 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2614 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2615 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2616 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2617 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2618 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2619 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2620 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2621 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2622 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2623 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2624 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2625 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2626 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2627 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2628 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2629 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2630 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2631 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R200 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M2632 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2633 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2634 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2635 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2636 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2637 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2638 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2639 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R201 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R202 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R203 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2640 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2641 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2642 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2643 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2644 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2645 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2646 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2647 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2648 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2649 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2650 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2651 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2652 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2653 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2654 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2655 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2656 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2657 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2658 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2659 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2660 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2661 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2662 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2663 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R204 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2664 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2665 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2666 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2667 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2668 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2669 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2670 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2671 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R205 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R206 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R207 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2672 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2673 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2674 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2675 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2676 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2677 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2678 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2679 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2680 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2681 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2682 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2683 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2684 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2685 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2686 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2687 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R208 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M2688 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2689 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2690 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2691 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2692 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2693 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2694 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2695 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R209 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R210 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R211 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2696 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2697 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2698 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2699 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2700 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2701 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2702 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2703 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2704 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2705 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2706 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2707 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2708 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2709 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2710 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2711 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2712 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2713 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2714 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2715 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2716 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2717 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2718 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2719 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R212 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2720 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2721 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2722 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2723 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2724 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2725 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2726 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2727 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R213 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R214 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R215 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2728 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2729 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2730 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2731 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2732 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2733 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2734 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2735 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2736 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2737 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2738 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2739 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2740 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2741 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2742 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2743 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2744 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2745 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2746 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2747 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2748 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2749 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2750 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2751 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R216 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M2752 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2753 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2754 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2755 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2756 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2757 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2758 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2759 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R217 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R218 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R219 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2760 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2761 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2762 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2763 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2764 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2765 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2766 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2767 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2768 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2769 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2770 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2771 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2772 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2773 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2774 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2775 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2776 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2777 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2778 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2779 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2780 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2781 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2782 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2783 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R220 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2784 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2785 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2786 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2787 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2788 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2789 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2790 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2791 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R221 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R222 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R223 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2792 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2793 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2794 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2795 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2796 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2797 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2798 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2799 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2800 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2801 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2802 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2803 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2804 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2805 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2806 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2807 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2808 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2809 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2810 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2811 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2812 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2813 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2814 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2815 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R224 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M2816 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2817 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2818 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2819 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2820 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2821 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2822 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2823 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R225 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R226 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R227 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2824 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2825 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2826 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2827 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2828 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2829 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2830 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2831 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2832 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2833 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2834 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2835 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2836 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2837 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2838 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2839 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2840 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2841 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2842 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2843 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2844 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2845 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2846 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2847 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R228 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2848 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2849 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2850 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2851 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2852 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2853 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2854 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2855 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R229 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R230 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R231 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2856 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2857 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2858 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2859 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2860 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2861 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2862 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2863 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2864 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2865 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2866 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2867 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2868 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2869 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2870 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2871 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2872 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2873 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2874 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2875 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2876 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2877 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2878 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2879 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R232 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M2880 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2881 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2882 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2883 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2884 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2885 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2886 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2887 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R233 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R234 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R235 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2888 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2889 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2890 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2891 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2892 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2893 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2894 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2895 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2896 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2897 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2898 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2899 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2900 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2901 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2902 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2903 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2904 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2905 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2906 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2907 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2908 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2909 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2910 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2911 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R236 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2912 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2913 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2914 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2915 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2916 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2917 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2918 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2919 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R237 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R238 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R239 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2920 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2921 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2922 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2923 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2924 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2925 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2926 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2927 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2928 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2929 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2930 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2931 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2932 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2933 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2934 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2935 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R240 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M2936 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2937 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2938 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2939 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2940 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2941 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2942 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2943 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R241 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R242 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R243 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2944 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2945 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2946 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2947 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2948 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2949 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2950 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2951 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2952 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2953 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2954 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2955 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2956 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2957 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2958 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2959 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2960 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2961 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2962 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2963 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2964 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2965 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2966 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2967 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R244 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2968 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2969 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2970 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2971 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2972 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2973 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2974 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2975 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R245 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R246 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R247 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2976 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2977 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2978 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2979 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2980 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2981 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2982 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2983 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2984 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2985 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2986 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2987 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2988 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2989 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2990 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2991 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2992 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2993 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2994 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2995 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2996 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2997 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2998 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2999 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R248 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M3000 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3001 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3002 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3003 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3004 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3005 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3006 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3007 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R249 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R250 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R251 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3008 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3009 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3010 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3011 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3012 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3013 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3014 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3015 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3016 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3017 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3018 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3019 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3020 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3021 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3022 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3023 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3024 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3025 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3026 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3027 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3028 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3029 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3030 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3031 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R252 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3032 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3033 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3034 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3035 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3036 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3037 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3038 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3039 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R253 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R254 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R255 8BitDac_1/R_in8 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3040 switchNew_0/a_86_24# D8 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3041 switchNew_0/a_105_21# switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3042 V_out9 switchNew_0/a_86_24# 8BitDac_0/V_out8 8BitDac_0/V_out8 pfet w=10 l=2
+  ad=140 pd=68 as=210 ps=102
M3043 8BitDac_0/V_out8 switchNew_0/a_105_21# V_out9 gnd nfet w=5 l=2
+  ad=137 pd=104 as=86 ps=64
M3044 switchNew_0/a_86_24# D8 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3045 switchNew_0/a_105_21# switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3046 V_out9 switchNew_0/a_86_24# 8BitDac_1/V_out8 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3047 V_out9 switchNew_0/a_105_21# 8BitDac_1/V_out8 V_out9 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3048 8BitDac_0/7BitDac_1/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3049 8BitDac_0/7BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3050 8BitDac_0/7BitDac_1/V_out7 8BitDac_0/7BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/V_out6 8BitDac_0/7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3051 8BitDac_0/7BitDac_1/6BitDac_0/V_out6 8BitDac_0/7BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/V_out7 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3052 8BitDac_0/7BitDac_1/switchNew_0/a_86_24# D6 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3053 8BitDac_0/7BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3054 8BitDac_0/7BitDac_1/V_out7 8BitDac_0/7BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3055 8BitDac_0/7BitDac_1/V_out7 8BitDac_0/7BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/V_out6 8BitDac_0/7BitDac_1/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3056 8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3057 8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3058 8BitDac_0/7BitDac_1/6BitDac_1/V_out6 8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3059 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3060 8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3061 8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3062 8BitDac_0/7BitDac_1/6BitDac_1/V_out6 8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3063 8BitDac_0/7BitDac_1/6BitDac_1/V_out6 8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 8BitDac_0/7BitDac_1/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3064 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3065 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3066 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3067 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3068 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3069 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3070 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3071 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3072 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3073 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3074 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3075 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3076 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3077 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3078 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3079 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3080 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3081 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3082 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3083 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3084 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3085 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3086 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_1/R_in8 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3087 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_1/R_in8 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R256 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_1/R_in8 polyResistor w=2 l=62
M3088 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3089 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3090 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3091 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3092 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3093 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3094 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3095 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R257 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R258 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R259 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3096 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3097 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3098 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3099 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3100 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3101 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3102 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3103 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3104 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3105 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3106 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3107 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3108 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3109 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3110 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3111 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3112 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3113 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3114 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3115 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3116 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3117 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3118 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3119 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R260 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3120 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3121 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3122 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3123 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3124 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3125 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3126 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3127 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R261 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R262 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R263 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3128 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3129 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3130 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3131 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3132 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3133 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3134 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3135 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3136 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3137 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3138 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3139 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3140 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3141 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3142 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3143 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3144 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3145 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3146 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3147 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3148 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3149 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3150 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3151 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R264 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M3152 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3153 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3154 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3155 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3156 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3157 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3158 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3159 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R265 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R266 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R267 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3160 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3161 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3162 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3163 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3164 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3165 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3166 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3167 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3168 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3169 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3170 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3171 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3172 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3173 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3174 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3175 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3176 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3177 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3178 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3179 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3180 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3181 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3182 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3183 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R268 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3184 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3185 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3186 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3187 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3188 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3189 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3190 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3191 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R269 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R270 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R271 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3192 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3193 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3194 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3195 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3196 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3197 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3198 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3199 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3200 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3201 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3202 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3203 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3204 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3205 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3206 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3207 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R272 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M3208 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3209 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3210 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3211 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3212 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3213 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3214 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3215 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R273 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R274 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R275 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3216 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3217 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3218 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3219 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3220 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3221 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3222 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3223 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3224 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3225 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3226 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3227 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3228 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3229 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3230 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3231 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3232 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3233 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3234 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3235 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3236 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3237 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3238 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3239 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R276 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3240 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3241 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3242 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3243 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3244 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3245 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3246 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3247 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R277 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R278 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R279 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3248 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3249 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3250 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3251 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3252 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3253 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3254 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3255 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3256 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3257 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3258 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3259 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3260 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3261 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3262 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3263 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3264 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3265 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3266 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3267 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3268 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3269 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3270 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3271 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R280 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M3272 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3273 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3274 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3275 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3276 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3277 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3278 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3279 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R281 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R282 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R283 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3280 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3281 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3282 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3283 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3284 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3285 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3286 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3287 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3288 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3289 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3290 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3291 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3292 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3293 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3294 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3295 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3296 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3297 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3298 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3299 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3300 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3301 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3302 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3303 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R284 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3304 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3305 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3306 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3307 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3308 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3309 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3310 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3311 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R285 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R286 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R287 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3312 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3313 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3314 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3315 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3316 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3317 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3318 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3319 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3320 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3321 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3322 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3323 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3324 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3325 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3326 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3327 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3328 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3329 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3330 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3331 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3332 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3333 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3334 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3335 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R288 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M3336 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3337 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3338 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3339 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3340 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3341 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3342 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3343 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R289 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R290 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R291 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3344 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3345 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3346 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3347 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3348 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3349 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3350 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3351 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3352 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3353 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3354 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3355 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3356 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3357 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3358 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3359 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3360 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3361 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3362 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3363 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3364 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3365 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3366 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3367 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R292 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3368 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3369 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3370 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3371 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3372 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3373 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3374 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3375 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R293 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R294 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R295 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3376 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3377 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3378 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3379 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3380 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3381 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3382 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3383 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3384 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3385 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3386 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3387 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3388 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3389 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3390 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3391 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3392 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3393 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3394 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3395 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3396 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3397 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3398 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3399 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R296 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M3400 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3401 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3402 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3403 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3404 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3405 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3406 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3407 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R297 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R298 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R299 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3408 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3409 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3410 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3411 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3412 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3413 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3414 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3415 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3416 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3417 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3418 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3419 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3420 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3421 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3422 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3423 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3424 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3425 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3426 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3427 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3428 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3429 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3430 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3431 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R300 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3432 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3433 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3434 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3435 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3436 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3437 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3438 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3439 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R301 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R302 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R303 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3440 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3441 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3442 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3443 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3444 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3445 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3446 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3447 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3448 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3449 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3450 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3451 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3452 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3453 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3454 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3455 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R304 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M3456 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3457 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3458 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3459 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3460 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3461 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3462 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3463 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R305 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R306 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R307 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3464 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3465 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3466 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3467 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3468 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3469 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3470 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3471 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3472 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3473 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3474 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3475 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3476 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3477 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3478 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3479 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3480 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3481 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3482 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3483 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3484 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3485 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3486 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3487 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R308 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3488 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3489 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3490 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3491 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3492 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3493 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3494 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3495 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R309 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R310 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R311 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3496 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3497 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3498 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3499 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3500 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3501 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3502 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3503 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3504 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3505 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3506 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3507 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3508 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3509 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3510 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3511 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3512 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3513 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3514 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3515 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3516 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3517 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3518 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3519 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R312 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M3520 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3521 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3522 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3523 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3524 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3525 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3526 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3527 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R313 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R314 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R315 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3528 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3529 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3530 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3531 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3532 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3533 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3534 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3535 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3536 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3537 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3538 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3539 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3540 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3541 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3542 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3543 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3544 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3545 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3546 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3547 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3548 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3549 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3550 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3551 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R316 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3552 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3553 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3554 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3555 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3556 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3557 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3558 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3559 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R317 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R318 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R319 8BitDac_0/7BitDac_1/6BitDac_1/R_in6 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3560 8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3561 8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3562 8BitDac_0/7BitDac_1/6BitDac_0/V_out6 8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3563 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3564 8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3565 8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3566 8BitDac_0/7BitDac_1/6BitDac_0/V_out6 8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3567 8BitDac_0/7BitDac_1/6BitDac_0/V_out6 8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 8BitDac_0/7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3568 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3569 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3570 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3571 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3572 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3573 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3574 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3575 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3576 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3577 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3578 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3579 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3580 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3581 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3582 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3583 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3584 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3585 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3586 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3587 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3588 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3589 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3590 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_1/R_in6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3591 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_1/R_in6 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R320 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_1/R_in6 polyResistor w=2 l=62
M3592 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3593 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3594 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3595 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3596 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3597 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3598 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3599 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R321 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R322 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R323 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3600 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3601 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3602 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3603 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3604 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3605 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3606 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3607 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3608 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3609 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3610 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3611 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3612 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3613 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3614 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3615 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3616 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3617 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3618 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3619 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3620 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3621 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3622 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3623 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R324 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3624 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3625 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3626 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3627 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3628 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3629 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3630 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3631 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R325 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R326 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R327 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3632 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3633 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3634 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3635 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3636 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3637 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3638 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3639 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3640 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3641 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3642 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3643 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3644 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3645 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3646 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3647 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3648 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3649 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3650 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3651 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3652 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3653 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3654 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3655 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R328 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M3656 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3657 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3658 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3659 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3660 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3661 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3662 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3663 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R329 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R330 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R331 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3664 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3665 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3666 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3667 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3668 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3669 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3670 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3671 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3672 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3673 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3674 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3675 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3676 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3677 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3678 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3679 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3680 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3681 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3682 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3683 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3684 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3685 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3686 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3687 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R332 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3688 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3689 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3690 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3691 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3692 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3693 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3694 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3695 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R333 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R334 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R335 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3696 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3697 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3698 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3699 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3700 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3701 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3702 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3703 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3704 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3705 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3706 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3707 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3708 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3709 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3710 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3711 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R336 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M3712 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3713 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3714 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3715 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3716 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3717 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3718 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3719 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R337 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R338 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R339 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3720 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3721 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3722 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3723 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3724 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3725 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3726 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3727 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3728 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3729 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3730 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3731 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3732 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3733 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3734 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3735 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3736 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3737 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3738 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3739 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3740 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3741 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3742 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3743 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R340 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3744 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3745 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3746 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3747 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3748 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3749 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3750 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3751 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R341 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R342 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R343 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3752 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3753 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3754 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3755 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3756 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3757 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3758 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3759 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3760 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3761 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3762 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3763 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3764 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3765 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3766 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3767 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3768 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3769 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3770 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3771 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3772 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3773 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3774 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3775 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R344 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M3776 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3777 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3778 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3779 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3780 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3781 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3782 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3783 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R345 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R346 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R347 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3784 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3785 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3786 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3787 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3788 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3789 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3790 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3791 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3792 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3793 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3794 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3795 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3796 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3797 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3798 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3799 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3800 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3801 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3802 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3803 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3804 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3805 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3806 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3807 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R348 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3808 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3809 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3810 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3811 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3812 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3813 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3814 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3815 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R349 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R350 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R351 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3816 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3817 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3818 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3819 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3820 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3821 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3822 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3823 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3824 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3825 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3826 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3827 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3828 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3829 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3830 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3831 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3832 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3833 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3834 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3835 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3836 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3837 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3838 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3839 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R352 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M3840 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3841 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3842 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3843 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3844 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3845 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3846 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3847 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R353 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R354 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R355 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3848 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3849 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3850 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3851 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3852 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3853 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3854 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3855 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3856 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3857 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3858 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3859 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3860 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3861 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3862 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3863 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3864 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3865 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3866 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3867 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3868 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3869 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3870 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3871 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R356 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3872 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3873 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3874 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3875 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3876 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3877 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3878 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3879 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R357 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R358 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R359 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3880 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3881 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3882 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3883 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3884 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3885 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3886 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3887 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3888 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3889 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3890 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3891 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3892 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3893 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3894 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3895 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3896 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3897 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3898 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3899 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3900 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3901 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3902 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3903 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R360 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M3904 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3905 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3906 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3907 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3908 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3909 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3910 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3911 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R361 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R362 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R363 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3912 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3913 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3914 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3915 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3916 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3917 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3918 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3919 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3920 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3921 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3922 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3923 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3924 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3925 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3926 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3927 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3928 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3929 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3930 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3931 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3932 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3933 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3934 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3935 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R364 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3936 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3937 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3938 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3939 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3940 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3941 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3942 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3943 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R365 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R366 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R367 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3944 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3945 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3946 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3947 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3948 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3949 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3950 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3951 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3952 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3953 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3954 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3955 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3956 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3957 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3958 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3959 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R368 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M3960 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3961 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3962 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3963 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3964 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3965 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3966 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3967 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R369 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R370 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R371 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3968 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3969 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3970 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3971 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3972 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3973 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3974 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3975 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3976 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3977 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3978 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3979 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3980 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3981 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3982 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3983 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3984 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3985 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3986 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3987 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3988 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3989 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3990 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3991 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R372 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3992 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3993 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3994 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3995 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3996 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3997 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3998 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3999 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R373 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R374 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R375 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4000 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4001 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4002 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4003 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4004 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4005 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4006 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4007 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4008 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4009 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4010 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4011 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4012 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4013 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4014 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4015 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4016 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4017 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4018 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4019 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4020 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4021 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4022 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4023 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R376 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M4024 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4025 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4026 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4027 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4028 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4029 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4030 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4031 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R377 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R378 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R379 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4032 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4033 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4034 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4035 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4036 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4037 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4038 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4039 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4040 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4041 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4042 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4043 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4044 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4045 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4046 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4047 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4048 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4049 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4050 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4051 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4052 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4053 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4054 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4055 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R380 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4056 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4057 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4058 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4059 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4060 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4061 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4062 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4063 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R381 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R382 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R383 8BitDac_0/7BitDac_1/R_in7 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4064 8BitDac_0/switchNew_0/a_86_24# D7 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4065 8BitDac_0/switchNew_0/a_105_21# 8BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4066 8BitDac_0/V_out8 8BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/V_out7 8BitDac_0/7BitDac_0/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4067 8BitDac_0/7BitDac_0/V_out7 8BitDac_0/switchNew_0/a_105_21# 8BitDac_0/V_out8 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4068 8BitDac_0/switchNew_0/a_86_24# D7 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4069 8BitDac_0/switchNew_0/a_105_21# 8BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4070 8BitDac_0/V_out8 8BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_1/V_out7 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4071 8BitDac_0/V_out8 8BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_1/V_out7 8BitDac_0/V_out8 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4072 8BitDac_0/7BitDac_0/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4073 8BitDac_0/7BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4074 8BitDac_0/7BitDac_0/V_out7 8BitDac_0/7BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/V_out6 8BitDac_0/7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4075 8BitDac_0/7BitDac_0/6BitDac_0/V_out6 8BitDac_0/7BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/V_out7 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4076 8BitDac_0/7BitDac_0/switchNew_0/a_86_24# D6 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4077 8BitDac_0/7BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4078 8BitDac_0/7BitDac_0/V_out7 8BitDac_0/7BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4079 8BitDac_0/7BitDac_0/V_out7 8BitDac_0/7BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/V_out6 8BitDac_0/7BitDac_0/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4080 8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4081 8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4082 8BitDac_0/7BitDac_0/6BitDac_1/V_out6 8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4083 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4084 8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4085 8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4086 8BitDac_0/7BitDac_0/6BitDac_1/V_out6 8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4087 8BitDac_0/7BitDac_0/6BitDac_1/V_out6 8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 8BitDac_0/7BitDac_0/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4088 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4089 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4090 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4091 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4092 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4093 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4094 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4095 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4096 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4097 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4098 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4099 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4100 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4101 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4102 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4103 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4104 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4105 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4106 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4107 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4108 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4109 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4110 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_1/R_in7 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4111 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_1/R_in7 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R384 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_1/R_in7 polyResistor w=2 l=62
M4112 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4113 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4114 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4115 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4116 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4117 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4118 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4119 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R385 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R386 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R387 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4120 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4121 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4122 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4123 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4124 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4125 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4126 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4127 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4128 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4129 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4130 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4131 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4132 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4133 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4134 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4135 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4136 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4137 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4138 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4139 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4140 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4141 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4142 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4143 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R388 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4144 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4145 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4146 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4147 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4148 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4149 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4150 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4151 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R389 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R390 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R391 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4152 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4153 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4154 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4155 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4156 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4157 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4158 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4159 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4160 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4161 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4162 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4163 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4164 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4165 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4166 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4167 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4168 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4169 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4170 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4171 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4172 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4173 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4174 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4175 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R392 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M4176 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4177 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4178 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4179 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4180 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4181 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4182 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4183 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R393 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R394 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R395 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4184 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4185 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4186 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4187 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4188 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4189 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4190 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4191 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4192 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4193 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4194 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4195 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4196 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4197 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4198 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4199 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4200 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4201 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4202 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4203 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4204 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4205 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4206 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4207 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R396 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4208 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4209 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4210 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4211 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4212 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4213 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4214 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4215 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R397 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R398 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R399 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4216 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4217 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4218 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4219 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4220 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4221 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4222 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4223 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4224 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4225 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4226 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4227 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4228 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4229 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4230 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4231 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R400 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M4232 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4233 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4234 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4235 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4236 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4237 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4238 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4239 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R401 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R402 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R403 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4240 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4241 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4242 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4243 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4244 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4245 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4246 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4247 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4248 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4249 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4250 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4251 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4252 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4253 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4254 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4255 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4256 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4257 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4258 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4259 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4260 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4261 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4262 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4263 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R404 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4264 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4265 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4266 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4267 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4268 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4269 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4270 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4271 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R405 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R406 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R407 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4272 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4273 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4274 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4275 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4276 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4277 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4278 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4279 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4280 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4281 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4282 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4283 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4284 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4285 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4286 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4287 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4288 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4289 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4290 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4291 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4292 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4293 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4294 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4295 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R408 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M4296 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4297 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4298 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4299 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4300 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4301 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4302 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4303 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R409 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R410 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R411 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4304 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4305 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4306 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4307 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4308 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4309 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4310 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4311 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4312 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4313 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4314 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4315 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4316 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4317 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4318 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4319 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4320 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4321 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4322 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4323 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4324 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4325 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4326 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4327 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R412 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4328 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4329 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4330 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4331 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4332 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4333 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4334 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4335 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R413 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R414 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R415 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4336 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4337 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4338 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4339 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4340 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4341 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4342 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4343 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4344 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4345 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4346 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4347 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4348 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4349 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4350 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4351 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4352 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4353 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4354 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4355 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4356 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4357 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4358 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4359 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R416 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M4360 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4361 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4362 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4363 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4364 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4365 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4366 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4367 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R417 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R418 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R419 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4368 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4369 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4370 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4371 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4372 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4373 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4374 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4375 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4376 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4377 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4378 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4379 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4380 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4381 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4382 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4383 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4384 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4385 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4386 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4387 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4388 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4389 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4390 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4391 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R420 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4392 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4393 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4394 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4395 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4396 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4397 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4398 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4399 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R421 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R422 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R423 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4400 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4401 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4402 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4403 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4404 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4405 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4406 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4407 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4408 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4409 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4410 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4411 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4412 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4413 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4414 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4415 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4416 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4417 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4418 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4419 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4420 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4421 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4422 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4423 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R424 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M4424 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4425 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4426 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4427 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4428 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4429 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4430 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4431 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R425 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R426 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R427 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4432 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4433 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4434 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4435 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4436 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4437 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4438 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4439 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4440 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4441 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4442 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4443 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4444 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4445 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4446 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4447 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4448 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4449 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4450 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4451 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4452 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4453 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4454 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4455 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R428 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4456 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4457 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4458 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4459 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4460 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4461 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4462 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4463 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R429 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R430 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R431 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4464 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4465 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4466 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4467 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4468 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4469 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4470 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4471 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4472 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4473 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4474 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4475 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4476 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4477 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4478 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4479 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R432 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M4480 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4481 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4482 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4483 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4484 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4485 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4486 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4487 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R433 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R434 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R435 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4488 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4489 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4490 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4491 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4492 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4493 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4494 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4495 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4496 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4497 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4498 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4499 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4500 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4501 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4502 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4503 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4504 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4505 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4506 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4507 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4508 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4509 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4510 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4511 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R436 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4512 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4513 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4514 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4515 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4516 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4517 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4518 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4519 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R437 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R438 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R439 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4520 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4521 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4522 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4523 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4524 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4525 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4526 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4527 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4528 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4529 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4530 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4531 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4532 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4533 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4534 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4535 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4536 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4537 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4538 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4539 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4540 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4541 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4542 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4543 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R440 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M4544 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4545 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4546 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4547 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4548 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4549 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4550 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4551 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R441 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R442 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R443 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4552 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4553 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4554 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4555 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4556 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4557 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4558 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4559 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4560 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4561 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4562 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4563 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4564 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4565 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4566 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4567 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4568 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4569 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4570 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4571 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4572 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4573 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4574 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4575 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R444 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4576 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4577 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4578 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4579 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4580 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4581 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4582 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4583 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R445 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R446 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R447 8BitDac_0/7BitDac_0/6BitDac_1/R_in6 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4584 8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4585 8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4586 8BitDac_0/7BitDac_0/6BitDac_0/V_out6 8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4587 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4588 8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4589 8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4590 8BitDac_0/7BitDac_0/6BitDac_0/V_out6 8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4591 8BitDac_0/7BitDac_0/6BitDac_0/V_out6 8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 8BitDac_0/7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4592 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4593 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4594 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4595 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4596 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4597 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4598 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4599 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4600 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4601 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4602 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4603 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4604 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4605 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4606 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4607 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4608 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4609 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4610 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4611 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4612 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4613 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4614 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_1/R_in6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4615 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_1/R_in6 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R448 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_1/R_in6 polyResistor w=2 l=62
M4616 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4617 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4618 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4619 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4620 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4621 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4622 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4623 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R449 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R450 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R451 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4624 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4625 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4626 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4627 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4628 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4629 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4630 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4631 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4632 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4633 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4634 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4635 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4636 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4637 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4638 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4639 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4640 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4641 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4642 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4643 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4644 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4645 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4646 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4647 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R452 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4648 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4649 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4650 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4651 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4652 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4653 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4654 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4655 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R453 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R454 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R455 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4656 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4657 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4658 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4659 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4660 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4661 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4662 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4663 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4664 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4665 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4666 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4667 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4668 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4669 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4670 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4671 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4672 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4673 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4674 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4675 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4676 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4677 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4678 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4679 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R456 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M4680 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4681 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4682 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4683 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4684 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4685 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4686 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4687 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R457 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R458 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R459 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4688 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4689 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4690 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4691 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4692 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4693 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4694 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4695 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4696 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4697 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4698 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4699 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4700 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4701 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4702 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4703 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4704 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4705 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4706 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4707 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4708 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4709 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4710 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4711 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R460 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4712 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4713 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4714 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4715 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4716 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4717 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4718 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4719 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R461 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R462 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R463 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4720 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4721 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4722 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4723 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4724 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4725 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4726 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4727 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4728 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4729 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4730 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4731 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4732 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4733 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4734 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4735 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R464 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M4736 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4737 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4738 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4739 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4740 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4741 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4742 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4743 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R465 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R466 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R467 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4744 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4745 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4746 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4747 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4748 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4749 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4750 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4751 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4752 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4753 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4754 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4755 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4756 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4757 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4758 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4759 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4760 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4761 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4762 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4763 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4764 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4765 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4766 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4767 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R468 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4768 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4769 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4770 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4771 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4772 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4773 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4774 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4775 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R469 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R470 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R471 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4776 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4777 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4778 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4779 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4780 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4781 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4782 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4783 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4784 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4785 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4786 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4787 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4788 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4789 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4790 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4791 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4792 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4793 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4794 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4795 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4796 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4797 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4798 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4799 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R472 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M4800 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4801 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4802 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4803 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4804 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4805 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4806 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4807 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R473 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R474 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R475 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4808 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4809 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4810 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4811 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4812 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4813 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4814 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4815 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4816 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4817 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4818 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4819 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4820 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4821 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4822 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4823 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4824 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4825 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4826 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4827 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4828 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4829 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4830 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4831 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R476 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4832 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4833 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4834 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4835 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4836 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4837 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4838 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4839 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R477 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R478 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R479 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4840 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4841 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4842 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4843 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4844 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4845 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4846 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4847 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4848 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4849 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4850 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4851 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4852 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4853 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4854 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4855 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4856 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4857 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4858 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4859 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4860 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4861 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4862 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4863 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R480 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M4864 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4865 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4866 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4867 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4868 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4869 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4870 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4871 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R481 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R482 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R483 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4872 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4873 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4874 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4875 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4876 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4877 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4878 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4879 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4880 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4881 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4882 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4883 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4884 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4885 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4886 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4887 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4888 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4889 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4890 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4891 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4892 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4893 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4894 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4895 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R484 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4896 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4897 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4898 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4899 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4900 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4901 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4902 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4903 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R485 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R486 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R487 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4904 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4905 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4906 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4907 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4908 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4909 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4910 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4911 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4912 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4913 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4914 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4915 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4916 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4917 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4918 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4919 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4920 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4921 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4922 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4923 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4924 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4925 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4926 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4927 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R488 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M4928 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4929 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4930 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4931 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4932 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4933 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4934 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4935 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R489 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R490 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R491 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4936 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4937 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4938 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4939 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4940 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4941 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4942 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4943 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4944 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4945 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4946 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4947 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4948 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4949 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4950 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4951 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4952 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4953 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4954 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4955 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4956 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4957 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4958 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4959 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R492 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4960 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4961 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4962 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4963 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4964 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4965 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4966 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4967 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R493 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R494 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R495 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4968 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4969 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4970 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4971 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4972 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4973 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4974 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4975 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4976 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4977 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4978 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4979 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4980 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4981 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4982 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4983 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R496 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M4984 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4985 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4986 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4987 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4988 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4989 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4990 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4991 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R497 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R498 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R499 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4992 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4993 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4994 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4995 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4996 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4997 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4998 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4999 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5000 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5001 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5002 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5003 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5004 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5005 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5006 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5007 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5008 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5009 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5010 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5011 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5012 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5013 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5014 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5015 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R500 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M5016 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5017 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5018 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5019 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5020 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5021 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5022 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5023 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R501 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R502 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R503 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M5024 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5025 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5026 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5027 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5028 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5029 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5030 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5031 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5032 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5033 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5034 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5035 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5036 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5037 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5038 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5039 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5040 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5041 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5042 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5043 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5044 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5045 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5046 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5047 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R504 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M5048 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5049 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5050 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5051 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5052 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5053 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5054 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5055 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R505 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R506 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R507 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M5056 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5057 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5058 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5059 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5060 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5061 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5062 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5063 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5064 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5065 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5066 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5067 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5068 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5069 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5070 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5071 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5072 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5073 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5074 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5075 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5076 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5077 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5078 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5079 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R508 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M5080 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5081 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5082 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5083 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5084 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5085 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5086 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5087 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R509 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R510 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R511 R_in9 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
C0 D6 8BitDac_0/7BitDac_0/6BitDac_0/V_out6 5.31fF
C1 D0 VA 20.85fF
C2 D2 VA 22.76fF
C3 D2 D1 116.51fF
C4 D2 8BitDac_0/7BitDac_0/V_out7 3.39fF
C5 D6 8BitDac_1/7BitDac_0/6BitDac_0/V_out6 5.31fF
C6 D6 8BitDac_0/7BitDac_1/6BitDac_0/V_out6 5.31fF
C7 D3 VA 31.46fF
C8 D3 D1 22.21fF
C9 D1 VA 61.14fF
C10 D4 VA 3.47fF
C11 D6 8BitDac_1/7BitDac_1/6BitDac_0/V_out6 5.31fF
C12 D5 gnd 2.49fF
C13 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C14 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C15 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C16 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C17 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C18 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C19 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C20 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C21 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C22 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C23 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C24 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C25 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C26 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C27 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C28 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C29 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C30 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C31 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C32 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C33 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C34 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C35 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C36 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C37 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C38 8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C39 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C40 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C41 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C42 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C43 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C44 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C45 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C46 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C47 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C48 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C49 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C50 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C51 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C52 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C53 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C54 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C55 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C56 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C57 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C58 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C59 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C60 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C61 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C62 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C63 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C64 8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C65 8BitDac_0/7BitDac_0/6BitDac_1/V_out6 gnd 2.06fF
C66 8BitDac_0/7BitDac_1/V_out7 gnd 2.40fF
C67 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C68 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C69 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C70 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C71 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C72 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C73 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C74 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C75 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C76 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C77 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C78 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C79 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C80 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C81 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C82 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C83 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C84 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C85 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C86 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C87 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C88 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C89 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C90 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C91 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C92 8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C93 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C94 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C95 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C96 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C97 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C98 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C99 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C100 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C101 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C102 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C103 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C104 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C105 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C106 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C107 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C108 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C109 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C110 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C111 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C112 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C113 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C114 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C115 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C116 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C117 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C118 8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C119 8BitDac_0/7BitDac_1/6BitDac_1/V_out6 gnd 2.06fF
C120 8BitDac_1/V_out8 gnd 2.32fF
C121 8BitDac_0/V_out8 gnd 2.04fF
C122 VA gnd 926.23fF
C123 8BitDac_1/R_in8 gnd 2.05fF
C124 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C125 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C126 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C127 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C128 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C129 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C130 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C131 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C132 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C133 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C134 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C135 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C136 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C137 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C138 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C139 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C140 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C141 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C142 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C143 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C144 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C145 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C146 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C147 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C148 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C149 8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C150 D1 gnd 77.30fF
C151 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C152 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C153 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C154 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C155 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C156 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C157 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C158 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C159 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C160 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C161 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C162 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C163 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C164 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C165 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C166 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C167 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C168 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C169 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C170 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C171 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C172 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C173 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C174 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C175 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C176 8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C177 8BitDac_1/7BitDac_0/6BitDac_1/V_out6 gnd 2.06fF
C178 8BitDac_1/7BitDac_1/V_out7 gnd 2.40fF
C179 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C180 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C181 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C182 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C183 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C184 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C185 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C186 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C187 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C188 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C189 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C190 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C191 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C192 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C193 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C194 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C195 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C196 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C197 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C198 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C199 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C200 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C201 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C202 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C203 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C204 8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C205 D0 gnd 101.47fF
C206 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C207 D2 gnd 61.63fF
C208 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C209 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C210 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C211 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C212 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C213 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C214 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C215 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C216 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C217 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C218 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C219 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C220 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C221 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C222 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C223 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C224 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C225 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C226 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C227 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C228 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C229 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C230 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C231 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C232 8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C233 8BitDac_1/7BitDac_1/6BitDac_1/V_out6 gnd 2.06fF




valpha  R_in9 Gnd 3.3
vbeta  VA Gnd 3.3
vzero D0 Gnd pulse(0 1.8 0.1m 60p 60p 0.1m 0.2m)
vone  D1 Gnd pulse(0 1.8 0.2m 60p 60p 0.2m 0.4m)
vtwo  D2 Gnd pulse(0 1.8 0.4m 60p 60p 0.4m 0.8m)
vthree D3 Gnd pulse(0 1.8 0.8m 60p 60p 0.8m 1.6m)
vfour D4 Gnd pulse (0 1.8 1.6m 60p 60p 1.6m 3.2m)
vfive D5 Gnd pulse (0 1.8 3.2m 60p 60p 3.2m 6.4m)
vsix D6 Gnd pulse (0 1.8 6.4m 60p 60p 6.4m 12.8m)
vseven D7 Gnd pulse (0 1.8 12.8m 60p 60p 12.8m 25.6m)
veight D8 Gnd pulse (0 1.8 25.6m 60p 60p 25.6m 51.2m)

.tran 0.01m 51.2m
.control
run

plot V(V_out9) V(D0)

.endc
.end






