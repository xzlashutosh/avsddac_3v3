magic
tech scmos
timestamp 1599308010
<< error_s >>
rect 2894 1619 2895 1620
<< metal1 >>
rect 16 3280 21 3283
rect 5 -23 11 -22
rect 5225 -23 5229 1
rect 5 -28 5229 -23
rect 5 -175 11 -28
rect 174 -119 177 -92
rect 1293 -147 1298 -57
rect 6146 -66 6149 1796
rect 6139 -102 6156 -98
rect 6266 -99 6302 -96
rect 6139 -132 6148 -129
rect 6139 -1630 6142 -132
rect 6280 -135 6283 -99
rect 6262 -139 6283 -135
rect 6262 -162 6274 -139
rect 6136 -1633 6142 -1630
rect 5214 -3427 5218 -3422
<< m2contact >>
rect 1293 -57 1298 -52
rect 174 -92 178 -85
rect 174 -126 178 -119
rect 1293 -152 1298 -147
<< metal2 >>
rect 2891 3385 2894 3387
rect 4399 3330 4419 3332
rect 4399 3328 4401 3330
rect 481 3292 484 3293
rect 1304 3273 1310 3280
rect 1974 3264 1977 3273
rect 6022 3227 6025 3230
rect 6010 1796 6025 1803
rect 6010 1672 6013 1796
rect 6010 1669 6119 1672
rect 480 1601 483 1623
rect 2882 1619 2895 1624
rect 480 1598 485 1601
rect 482 -133 485 1598
rect 2882 1537 2887 1619
rect 2882 1532 2974 1537
rect 1293 1402 1309 1406
rect 1293 -52 1298 1402
rect 2969 1291 2974 1532
rect 2845 1286 2974 1291
rect 2845 -39 2850 1286
rect 6116 1281 6119 1669
rect 6011 1278 6119 1281
rect 2880 -39 2885 -38
rect 2845 -42 2886 -39
rect 2880 -43 2885 -42
rect 470 -136 485 -133
rect 1293 -147 1298 -146
rect 6011 -199 6014 1278
<< m3contact >>
rect 174 -92 178 -85
rect 174 -126 178 -119
rect 1293 -152 1298 -147
<< metal3 >>
rect 344 3353 350 3356
rect 981 3347 989 3351
rect 175 3319 179 3323
rect 1585 3313 1589 3318
rect 184 3304 185 3307
rect 1678 3282 1681 3286
rect 40 3271 44 3274
rect 1533 3255 1537 3257
rect 690 3245 694 3252
rect 824 3202 825 3209
rect 836 3205 841 3210
rect 326 735 330 833
rect 326 731 470 735
rect 167 232 174 235
rect 167 228 170 232
rect 171 228 174 232
rect 167 225 291 228
rect 288 202 291 225
rect 288 199 385 202
rect 27 82 31 95
rect 27 78 33 82
rect 29 -155 33 78
rect 162 -106 166 132
rect 382 52 385 199
rect 174 49 385 52
rect 174 -85 177 49
rect 333 -73 339 -71
rect 466 -89 470 731
rect 162 -107 168 -106
rect 162 -109 166 -107
<< metal4 >>
rect 163 3337 171 3339
rect 1644 3329 1648 3331
rect 810 3238 815 3241
rect 1655 3233 1661 3236
rect 161 380 164 430
rect 158 377 164 380
rect 158 -66 161 377
rect 153 -74 161 -66
rect 152 -84 161 -74
rect 152 -89 160 -84
<< metal5 >>
rect 115 3227 122 3239
rect 1608 3210 1615 3217
rect 6090 -51 6182 -46
rect 104 -197 111 -191
rect 6090 -253 6095 -51
rect 6177 -61 6182 -51
rect 5401 -258 6095 -253
<< metal6 >>
rect 6168 -142 6175 -136
rect 6168 -1723 6174 -142
rect 6085 -1729 6174 -1723
rect 5255 -3447 5260 -3428
use 9BitDac  9BitDac_0
timestamp 1599295951
transform 1 0 0 0 1 7
box 0 -40 6147 3379
use 9BitDac  9BitDac_1
timestamp 1599295951
transform 1 0 -11 0 1 -3419
box 0 -40 6147 3379
use switchNew  switchNew_0
timestamp 1599222484
transform 1 0 6079 0 1 -138
box 69 -1 187 81
use capacitor2  capacitor2_0
timestamp 1599096684
transform 0 1 6162 -1 0 -267
box -105 -12 219 150
<< labels >>
rlabel metal1 5214 -3427 5218 -3427 1 gnd!
rlabel metal1 16 3282 21 3282 1 R_in10
rlabel metal1 6150 -102 6150 -98 1 D9!
rlabel metal1 6302 -99 6302 -96 7 V_out10
rlabel metal6 5255 -3447 5260 -3447 1 gnd
rlabel metal4 163 3339 171 3339 1 D3
rlabel metal3 175 3322 179 3322 1 D1
rlabel metal3 184 3304 184 3307 1 D2
rlabel metal5 115 3229 122 3229 1 VA
rlabel metal3 344 3356 350 3356 1 D4
rlabel metal2 481 3293 484 3293 1 D5
rlabel metal2 1304 3280 1310 3280 1 D6
rlabel metal2 2891 3387 2894 3387 5 D7
rlabel metal2 6022 3230 6025 3230 1 D8
rlabel metal3 29 -151 33 -151 1 D0
rlabel metal4 152 -87 160 -87 1 D3
rlabel metal3 164 -106 168 -106 1 D1
rlabel metal3 333 -71 339 -71 1 D4
rlabel metal2 470 -133 473 -133 1 D5
rlabel metal2 1293 -146 1298 -146 1 D6
rlabel metal2 2880 -38 2885 -38 1 D7
rlabel metal2 6011 -196 6014 -196 1 D8
rlabel metal5 104 -197 111 -197 1 VA!
rlabel metal5 115 3227 122 3227 1 VA!
rlabel metal3 40 3274 44 3274 1 D0!
rlabel metal3 175 3323 179 3323 1 D1!
rlabel metal3 690 3252 694 3252 1 D0!
rlabel metal4 810 3238 810 3241 1 D3!
rlabel metal3 824 3202 824 3209 1 D1!
rlabel metal3 841 3205 841 3210 1 D2!
rlabel metal3 981 3351 989 3351 1 D4!
rlabel metal3 1533 3257 1537 3257 1 D0!
rlabel metal5 1608 3210 1615 3210 1 VA
rlabel metal4 1661 3233 1661 3236 1 D3
rlabel metal3 1585 3318 1589 3318 1 D1
rlabel metal4 1644 3331 1648 3331 1 D3
rlabel metal3 1678 3286 1681 3286 1 D2
rlabel space 1974 3272 1978 3272 1 D5
<< end >>
