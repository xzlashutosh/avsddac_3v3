* SPICE3 file created from 7BitDac.ext - technology: scmos
.model polyResistor R ( TC1=0 TC2=0 RSH=7.7 DEFW=1.E-7 NARROW=0.0 TNOM=27)

.model pfet PMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=4.1589E17 VTH0=-0.3938813 K1=0.5479015 K2=0.0360586 K3=0.0993095 K3B=5.7086622 W0=1E-6 NLX=1.313191E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=0.4911363 DVT1=0.2227356 DVT2=0.1 U0=115.6852975 UA=1.505832E-9 UB=1E-21 UC=-1E-10 VSAT=1.329694E5 A0=1.7590478 AGS=0.3641621 B0=3.427126E-7 B1=1.062928E-6 KETA=0.0134667 A1=0.6859506 A2=0.3506788 RDSW=168.5705677 PRWG=0.5 PRWB=-0.4987371 WR=1 WINT=0 LINT=3.028832E-8 XL=0 XW=-1E-8 DWG=-2.349633E-8 DWB=-7.152486E-9 VOFF=-0.0994037 NFACTOR=1.9424315 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=0.0608072 ETAB=-0.0426148 DSUB=0.7343015 PCLM=3.2579974 PDIBLC1=7.229527E-6 PDIBLC2=0.025389 PDIBLCB=-1E-3 DROUT=0 PSCBE1=1.454878E10 PSCBE2=4.202027E-9 PVAG=15 DELTA=0.01 RSH=7.8 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=6.32E-10 CGSO=6.32E-10 CGBO=1E-12 CJ=1.172138E-3 PB=0.8421173 MJ=0.4109788 CJSW=2.242609E-10 PBSW=0.8 MJSW=0.3752089 CJSWG=4.22E-10 PBSWG=0.8 MJSWG=0.3752089 CF=0 PVTH0=1.888482E-3 PRDSW=11.5315407 PK2=1.559399E-3 WKETA=0.0319301 LKETA=2.955547E-3 PU0=-1.1105313 PUA=-4.62102E-11 PUB=1E-21 PVSAT=50 PETA0=1E-4 PKETA=-4.346368E-3)

.model nfet NMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=2.3549E17 VTH0=0.3823463 K1=0.5810697 K2=4.774618E-3 K3=0.0431669 K3B=1.1498346 W0=1E-7 NLX=1.910552E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=1.2894824 DVT1=0.3622063 DVT2=0.0713729 U0=280.633249 UA=-1.208537E-9 UB=2.158625E-18 UC=5.342807E-11 VSAT=9.366802E4 A0=1.7593146 AGS=0.3939741 B0=-6.413949E-9 B1=-1E-7 KETA=-5.180424E-4 A1=0 A2=1 RDSW=105.5517558 PRWG=0.5 PRWB=-0.1998871 WR=1 WINT=7.904732E-10 LINT=1.571424E-8 XL=0 XW=-1E-8 DWG=1.297221E-9 DWB=1.479041E-9 VOFF=-0.0955434 NFACTOR=2.4358891 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=3.104851E-3 ETAB=-2.512384E-5 DSUB=0.0167075 PCLM=0.8073191 PDIBLC1=0.1666161 PDIBLC2=3.112892E-3 PDIBLCB=-0.1 DROUT=0.7875618 PSCBE1=8E10 PSCBE2=9.213635E-10 PVAG=3.85243E-3 DELTA=0.01 RSH=6.7 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=7.08E-10 CGSO=7.08E-10 CGBO=1E-12 CJ=9.68858E-4 PB=0.8 MJ=0.3864502 CJSW=2.512138E-10 PBSW=0.809286 MJSW=0.1060414 CJSWG=3.3E-10 PBSWG=0.809286 MJSWG=0.1060414 CF=0 PVTH0=-1.192722E-3 PRDSW=-5 PK2=6.450505E-5 WKETA=-4.27294E-4 LKETA=-0.0104078 PU0=6.3268729 PUA=2.226552E-11 PUB=0 PVSAT=969.1480157 PETA0=1E-4 PKETA=-1.049509E-3)


.option scale=0.1u

M1000 switchNew_0/a_86_24# D6 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=17780 ps=8636
M1001 switchNew_0/a_105_20# switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1002 V_out7 switchNew_0/a_86_24# 6BitDac_0/V_out6 6BitDac_0/V_out6 pfet w=10 l=2
+  ad=140 pd=68 as=210 ps=102
M1003 6BitDac_0/V_out6 switchNew_0/a_105_20# V_out7 gnd nfet w=5 l=2
+  ad=137 pd=104 as=86 ps=64
M1004 switchNew_0/a_86_24# D6 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=8890 ps=6096
M1005 switchNew_0/a_105_20# switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1006 V_out7 switchNew_0/a_86_24# 6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1007 V_out7 switchNew_0/a_105_20# 6BitDac_1/V_out6 V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1008 6BitDac_1/switchNew_0/a_86_24# D5 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1009 6BitDac_1/switchNew_0/a_105_20# 6BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1010 6BitDac_1/V_out6 6BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/V_out5 6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1011 6BitDac_1/5BitDac_0/V_out5 6BitDac_1/switchNew_0/a_105_20# 6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1012 6BitDac_1/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1013 6BitDac_1/switchNew_0/a_105_20# 6BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1014 6BitDac_1/V_out6 6BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1015 6BitDac_1/V_out6 6BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/V_out5 6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1016 6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1017 6BitDac_1/5BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1018 6BitDac_1/5BitDac_1/V_out5 6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/V_out4 6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1019 6BitDac_1/5BitDac_1/4BitDac_0/V_out4 6BitDac_1/5BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1020 6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1021 6BitDac_1/5BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1022 6BitDac_1/5BitDac_1/V_out5 6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1023 6BitDac_1/5BitDac_1/V_out5 6BitDac_1/5BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/V_out4 6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1024 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1025 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1026 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1027 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1028 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1029 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1030 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1031 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1032 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1033 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1034 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1035 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1036 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1037 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1038 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# R_out7 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1039 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# R_out7 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R0 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma R_out7 polyResistor w=2 l=62
R1 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
M1040 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1041 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1042 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1043 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1044 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1045 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1046 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1047 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R3 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1048 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1049 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1050 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1051 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1052 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1053 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1054 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1055 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1056 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1057 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1058 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1059 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1060 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1061 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1062 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1063 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1064 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1065 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1066 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1067 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1068 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1069 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1070 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1071 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R4 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
R5 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
M1072 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1073 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1074 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1075 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1076 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1077 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1078 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1079 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R6 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R7 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1080 6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1081 6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1082 6BitDac_1/5BitDac_1/4BitDac_1/V_out4 6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1083 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1084 6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1085 6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1086 6BitDac_1/5BitDac_1/4BitDac_1/V_out4 6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 6BitDac_1/5BitDac_1/4BitDac_1/V_out4 6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1089 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1090 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1091 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1092 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1093 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1094 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1095 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1096 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1097 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1098 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1099 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1100 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1101 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1102 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1103 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R8 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
R9 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
M1104 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1105 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1106 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1107 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1108 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1109 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1110 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1111 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R10 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R11 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1112 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1113 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1114 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1115 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1116 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1117 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1118 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1120 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1121 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1122 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1123 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1124 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1125 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1126 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1127 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1128 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1129 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1130 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1131 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1132 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1133 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1134 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1135 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R12 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
R13 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
M1136 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1137 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1138 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1139 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1140 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1141 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1142 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1143 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R14 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R15 6BitDac_1/5BitDac_1/4BitDac_1/R_in4 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1144 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1145 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1146 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1147 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1148 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1149 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1150 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1151 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1152 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1153 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1154 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1155 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1156 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1157 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1158 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1159 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_1/R_in4 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R16 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
R17 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
M1160 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1161 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1162 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1163 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1164 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1165 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1166 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1167 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R18 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R19 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1168 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1169 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1170 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1171 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1172 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1173 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1174 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1177 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1178 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1179 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1180 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1181 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1182 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1183 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1184 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1185 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1186 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1187 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1188 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1189 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1190 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1191 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R20 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
R21 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
M1192 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1193 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1194 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1195 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1196 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1197 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1198 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1199 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R22 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R23 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1200 6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1201 6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1202 6BitDac_1/5BitDac_1/4BitDac_0/V_out4 6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1203 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1204 6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1205 6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1206 6BitDac_1/5BitDac_1/4BitDac_0/V_out4 6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 6BitDac_1/5BitDac_1/4BitDac_0/V_out4 6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1209 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1210 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1211 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1212 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1213 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1214 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1215 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1216 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1217 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1218 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1219 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1220 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1221 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1222 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1223 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R24 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
R25 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
M1224 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1225 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1226 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1227 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1228 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1229 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1230 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1231 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R26 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R27 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1232 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1233 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1234 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1235 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1236 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1237 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1238 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1240 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1241 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1242 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1243 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1244 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1245 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1246 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1247 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1248 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1249 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1250 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1251 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1252 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1253 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1254 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1255 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R28 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
R29 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
M1256 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1257 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1258 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1259 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1260 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1261 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1262 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1263 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R30 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R31 6BitDac_1/5BitDac_1/R_in5 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1264 6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1265 6BitDac_1/5BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1266 6BitDac_1/5BitDac_0/V_out5 6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/V_out4 6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1267 6BitDac_1/5BitDac_0/4BitDac_0/V_out4 6BitDac_1/5BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1268 6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1269 6BitDac_1/5BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1270 6BitDac_1/5BitDac_0/V_out5 6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1271 6BitDac_1/5BitDac_0/V_out5 6BitDac_1/5BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/V_out4 6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1272 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1273 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1274 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1275 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1276 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1277 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1278 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1279 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1280 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1281 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1282 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1283 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1284 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1285 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1286 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1287 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_1/R_in5 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R32 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
R33 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
M1288 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1289 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1290 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1291 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1292 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1293 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1294 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1295 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R34 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R35 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1296 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1297 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1298 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1299 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1300 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1301 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1302 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1303 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1304 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1305 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1306 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1307 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1308 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1309 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1310 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1311 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1312 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1313 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1314 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1315 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1316 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1317 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1318 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1319 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R36 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
R37 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
M1320 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1321 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1322 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1323 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1324 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1325 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1326 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1327 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R38 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R39 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1328 6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1329 6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1330 6BitDac_1/5BitDac_0/4BitDac_1/V_out4 6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1331 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1332 6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1333 6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1334 6BitDac_1/5BitDac_0/4BitDac_1/V_out4 6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1335 6BitDac_1/5BitDac_0/4BitDac_1/V_out4 6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1336 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1337 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1338 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1339 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1340 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1341 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1342 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1343 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1344 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1345 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1346 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1347 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1348 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1349 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1350 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1351 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R40 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
R41 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
M1352 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1353 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1354 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1355 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1356 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1357 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1358 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1359 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R42 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R43 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1360 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1361 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1362 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1363 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1364 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1365 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1366 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1367 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1368 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1369 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1370 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1371 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1372 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1373 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1374 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1375 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1376 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1377 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1378 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1379 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1380 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1381 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1382 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1383 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R44 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
R45 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
M1384 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1385 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1386 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1387 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1388 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1389 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1390 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1391 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R46 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R47 6BitDac_1/5BitDac_0/4BitDac_1/R_in4 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1392 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1393 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1394 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1395 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1396 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1397 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1398 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1399 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1400 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1401 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1402 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1403 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1404 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1405 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1406 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1407 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_1/R_in4 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R48 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
R49 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
M1408 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1409 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1410 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1411 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1412 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1413 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1414 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1415 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R50 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R51 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1416 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1417 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1418 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1419 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1420 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1421 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1422 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1423 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1424 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1425 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1426 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1427 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1428 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1429 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1430 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1431 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1432 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1433 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1434 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1435 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1436 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1437 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1438 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1439 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R52 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
R53 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
M1440 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1441 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1442 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1443 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1444 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1445 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1446 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1447 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R54 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R55 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1448 6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1449 6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1450 6BitDac_1/5BitDac_0/4BitDac_0/V_out4 6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1451 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1452 6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1453 6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1454 6BitDac_1/5BitDac_0/4BitDac_0/V_out4 6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1455 6BitDac_1/5BitDac_0/4BitDac_0/V_out4 6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1456 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1457 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1458 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1459 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1460 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1461 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1462 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1463 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1464 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1465 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1466 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1467 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1468 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1469 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1470 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1471 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R56 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
R57 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
M1472 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1473 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1474 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1475 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1476 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1477 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1478 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1479 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R58 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R59 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1480 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1481 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1482 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1483 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1484 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1485 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1486 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1487 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1488 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1489 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1490 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1491 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1492 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1493 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1494 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1495 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1496 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1497 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1498 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1499 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1500 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1501 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1502 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1503 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R60 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
R61 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
M1504 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1505 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1506 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1507 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1508 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1509 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1510 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1511 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R62 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R63 6BitDac_1/R_in6 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1512 6BitDac_0/switchNew_0/a_86_24# D5 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1513 6BitDac_0/switchNew_0/a_105_20# 6BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1514 6BitDac_0/V_out6 6BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/V_out5 6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1515 6BitDac_0/5BitDac_0/V_out5 6BitDac_0/switchNew_0/a_105_20# 6BitDac_0/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1516 6BitDac_0/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1517 6BitDac_0/switchNew_0/a_105_20# 6BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1518 6BitDac_0/V_out6 6BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1519 6BitDac_0/V_out6 6BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/V_out5 6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1520 6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1521 6BitDac_0/5BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1522 6BitDac_0/5BitDac_1/V_out5 6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/V_out4 6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1523 6BitDac_0/5BitDac_1/4BitDac_0/V_out4 6BitDac_0/5BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1524 6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1525 6BitDac_0/5BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1526 6BitDac_0/5BitDac_1/V_out5 6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1527 6BitDac_0/5BitDac_1/V_out5 6BitDac_0/5BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/V_out4 6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1528 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1529 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1530 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1531 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1532 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1533 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1534 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1535 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1536 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1537 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1538 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1539 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1540 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1541 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1542 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_1/R_in6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1543 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_1/R_in6 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R64 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 6BitDac_1/R_in6 polyResistor w=2 l=62
R65 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
M1544 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1545 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1546 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1547 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1548 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1549 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1550 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1551 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R66 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R67 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1552 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1553 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1554 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1555 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1556 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1557 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1558 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1559 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1560 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1561 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1562 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1563 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1564 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1565 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1566 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1567 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1568 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1569 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1570 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1571 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1572 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1573 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1574 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1575 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R68 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
R69 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
M1576 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1577 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1578 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1579 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1580 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1581 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1582 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1583 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R70 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R71 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1584 6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1585 6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1586 6BitDac_0/5BitDac_1/4BitDac_1/V_out4 6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1587 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1588 6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1589 6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1590 6BitDac_0/5BitDac_1/4BitDac_1/V_out4 6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1591 6BitDac_0/5BitDac_1/4BitDac_1/V_out4 6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1592 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1593 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1594 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1595 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1596 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1597 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1598 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1599 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1600 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1601 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1602 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1603 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1604 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1605 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1606 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1607 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R72 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
R73 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
M1608 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1609 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1610 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1611 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1612 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1613 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1614 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1615 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R74 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R75 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1616 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1617 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1618 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1619 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1620 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1621 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1622 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1623 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1624 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1625 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1626 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1627 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1628 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1629 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1630 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1631 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1632 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1633 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1634 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1635 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1636 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1637 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1638 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1639 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R76 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
R77 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
M1640 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1641 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1642 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1643 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1644 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1645 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1646 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1647 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R78 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R79 6BitDac_0/5BitDac_1/4BitDac_1/R_in4 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1648 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1649 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1650 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1651 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1652 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1653 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1654 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1655 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1656 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1657 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1658 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1659 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1660 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1661 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1662 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1663 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_1/R_in4 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R80 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
R81 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
M1664 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1665 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1666 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1667 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1668 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1669 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1670 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1671 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R82 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R83 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1672 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1673 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1674 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1675 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1676 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1677 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1678 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1679 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1680 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1681 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1682 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1683 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1684 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1685 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1686 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1687 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1688 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1689 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1690 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1691 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1692 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1693 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1694 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1695 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R84 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
R85 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
M1696 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1697 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1698 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1699 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1700 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1701 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1702 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1703 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R86 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R87 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1704 6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1705 6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1706 6BitDac_0/5BitDac_1/4BitDac_0/V_out4 6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1707 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1708 6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1709 6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1710 6BitDac_0/5BitDac_1/4BitDac_0/V_out4 6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1711 6BitDac_0/5BitDac_1/4BitDac_0/V_out4 6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1712 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1713 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1714 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1715 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1716 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1717 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1718 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1719 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1720 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1721 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1722 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1723 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1724 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1725 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1726 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1727 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R88 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
R89 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
M1728 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1729 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1730 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1731 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1732 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1733 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1734 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1735 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R90 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R91 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1736 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1737 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1738 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1739 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1740 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1741 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1742 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1743 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1744 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1745 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1746 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1747 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1748 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1749 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1750 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1751 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1752 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1753 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1754 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1755 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1756 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1757 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1758 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1759 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R92 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
R93 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
M1760 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1761 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1762 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1763 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1764 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1765 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1766 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1767 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R94 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R95 6BitDac_0/5BitDac_1/R_in5 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1768 6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1769 6BitDac_0/5BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1770 6BitDac_0/5BitDac_0/V_out5 6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/V_out4 6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1771 6BitDac_0/5BitDac_0/4BitDac_0/V_out4 6BitDac_0/5BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1772 6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1773 6BitDac_0/5BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1774 6BitDac_0/5BitDac_0/V_out5 6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1775 6BitDac_0/5BitDac_0/V_out5 6BitDac_0/5BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/V_out4 6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1776 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1777 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1778 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1779 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1780 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1781 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1782 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1783 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1784 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1785 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1786 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1787 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1788 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1789 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1790 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1791 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_1/R_in5 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R96 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
R97 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
M1792 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1793 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1794 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1795 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1796 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1797 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1798 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1799 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R98 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R99 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1800 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1801 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1802 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1803 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1804 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1805 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1806 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1807 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1808 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1809 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1810 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1811 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1812 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1813 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1814 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1815 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1816 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1817 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1818 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1819 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1820 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1821 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1822 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1823 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R100 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
R101 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
M1824 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1825 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1826 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1827 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1828 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1829 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1830 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1831 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R102 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R103 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1832 6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1833 6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1834 6BitDac_0/5BitDac_0/4BitDac_1/V_out4 6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1835 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1836 6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1837 6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1838 6BitDac_0/5BitDac_0/4BitDac_1/V_out4 6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1839 6BitDac_0/5BitDac_0/4BitDac_1/V_out4 6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1840 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1841 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1842 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1843 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1844 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1845 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1846 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1847 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1848 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1849 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1850 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1851 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1852 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1853 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1854 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1855 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R104 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
R105 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
M1856 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1857 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1858 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1859 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1860 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1861 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1862 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1863 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R106 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R107 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1864 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1865 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1866 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1867 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1868 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1869 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1870 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1871 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1872 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1873 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1874 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1875 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1876 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1877 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1878 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1879 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1880 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1881 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1882 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1883 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1884 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1885 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1886 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1887 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R108 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
R109 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
M1888 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1889 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1890 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1891 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1892 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1893 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1894 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1895 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R110 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R111 6BitDac_0/5BitDac_0/4BitDac_1/R_in4 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1896 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1897 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1898 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1899 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1900 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1901 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1902 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1903 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1904 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1905 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1906 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1907 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1908 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1909 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1910 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1911 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_1/R_in4 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R112 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
R113 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
M1912 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1913 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1914 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1915 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1916 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1917 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1918 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1919 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R114 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R115 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1920 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1921 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1922 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1923 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1924 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1925 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1926 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1927 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1928 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1929 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1930 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1931 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1932 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1933 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1934 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1935 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1936 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1937 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1938 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1939 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1940 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1941 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1942 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1943 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R116 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
R117 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
M1944 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1945 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1946 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1947 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1948 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1949 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1950 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1951 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R118 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R119 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1952 6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1953 6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1954 6BitDac_0/5BitDac_0/4BitDac_0/V_out4 6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1955 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1956 6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1957 6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1958 6BitDac_0/5BitDac_0/4BitDac_0/V_out4 6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1959 6BitDac_0/5BitDac_0/4BitDac_0/V_out4 6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1960 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1961 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1962 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1963 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1964 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1965 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1966 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1967 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1968 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1969 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1970 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1971 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1972 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1973 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1974 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1975 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R120 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
R121 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
M1976 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1977 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1978 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1979 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1980 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1981 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1982 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1983 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R122 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R123 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1984 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1985 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1986 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1987 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1988 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1989 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1990 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1991 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1992 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1993 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1994 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1995 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1996 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1997 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1998 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1999 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2000 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2001 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2002 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2003 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2004 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2005 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2006 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2007 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R124 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
R125 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
M2008 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2009 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# Vdd Vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2010 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2011 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2012 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2013 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2014 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2015 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_20# 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R126 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R127 R_in7 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
C0 D1 D3 11.94fF
C1 D6 6BitDac_0/V_out6 5.31fF
C2 Vdd D2 2.71fF
C3 Vdd D0 4.30fF
C4 D2 D1 30.57fF
C5 Vdd D1 2.52fF
C6 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.17fF
C7 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C8 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C9 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.22fF
C10 6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd 2.30fF
C11 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.17fF
C12 6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C13 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.17fF
C14 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C15 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C16 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.22fF
C17 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.17fF
C18 6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C19 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.17fF
C20 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C21 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C22 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.22fF
C23 6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd 2.30fF
C24 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.17fF
C25 6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C26 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.17fF
C27 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C28 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C29 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.22fF
C30 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.17fF
C31 6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C32 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.17fF
C33 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C34 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C35 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.22fF
C36 6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd 2.30fF
C37 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.17fF
C38 6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C39 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.17fF
C40 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C41 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C42 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.22fF
C43 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.17fF
C44 6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C45 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.17fF
C46 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C47 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C48 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.22fF
C49 D3 gnd 2.24fF
C50 6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd 2.30fF
C51 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.17fF
C52 6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C53 D1 gnd 12.50fF
C54 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.17fF
C55 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C56 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C57 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.22fF
C58 D0 gnd 20.37fF
C59 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.17fF
C60 D2 gnd 5.32fF
C61 6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C62 D4 gnd 4.02fF
C63 6BitDac_1/V_out6 gnd 2.07fF
C64 Vdd gnd 122.48fF

valpha  R_in7 R_out7 3.3
vbeta  Vdd Gnd 3.3
vzero D0 Gnd pulse(0 1.8 0.1m 60p 60p 0.1m 0.2m)
vone  D1 Gnd pulse(0 1.8 0.2m 60p 60p 0.2m 0.4m)
vtwo  D2 Gnd pulse(0 1.8 0.4m 60p 60p 0.4m 0.8m)
vthree D3 Gnd pulse(0 1.8 0.8m 60p 60p 0.8m 1.6m)
vfour D4 Gnd pulse (0 1.8 1.6m 60p 60p 1.6m 3.2m)
vfive D5 Gnd pulse (0 1.8 3.2m 60p 60p 3.2m 6.4m)
vsix D6 Gnd pulse (0 1.8 6.4m 60p 60p 6.4m 12.8m)

.tran 0.01m 12.8m
.control
run

plot V(V_out7) V(D0)

.endc
.end

