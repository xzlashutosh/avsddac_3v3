magic
tech scmos
timestamp 1599268620
<< metal1 >>
rect 1429 3326 2890 3329
rect 968 3286 1000 3289
rect 969 3273 1001 3276
rect 1351 3256 1362 3259
rect 16 3241 21 3249
rect 709 3219 1268 3224
rect 1429 1381 1433 3326
rect 1686 3248 1692 3253
rect 1624 3242 1692 3248
rect 1412 1378 1433 1381
rect 1429 1377 1433 1378
rect 1487 3221 1514 3224
rect 1487 2 1491 3221
rect 2887 1625 2890 3326
rect 2887 1622 2898 1625
rect 2896 1586 2906 1590
rect 3016 1589 3020 1592
rect 2892 1556 2898 1559
rect 2892 1460 2895 1556
rect 2892 1457 2931 1460
rect 2928 1362 2931 1457
rect 2925 1359 2931 1362
rect 669 -1 1491 2
rect 2162 -20 2166 -18
<< m2contact >>
rect 961 3286 968 3290
rect 1000 3284 1007 3292
rect 962 3273 969 3277
rect 1001 3272 1008 3280
rect 1347 3256 1351 3260
rect 1362 3256 1366 3260
rect 705 3219 709 3224
rect 1268 3219 1273 3224
rect 1686 3253 1692 3258
rect 1615 3237 1624 3249
rect 2891 1586 2896 1590
<< metal2 >>
rect 1355 3308 2801 3311
rect 481 3258 484 3262
rect 1130 3256 1347 3259
rect 1304 3249 1309 3251
rect 1355 3249 1358 3308
rect 1366 3256 1634 3259
rect 1304 3245 1358 3249
rect 1631 3239 1634 3256
rect 1631 3236 1976 3239
rect 1631 3235 1634 3236
rect 2797 3230 2801 3308
rect 2891 1590 2894 3332
<< m3contact >>
rect 961 3286 968 3290
rect 1000 3284 1007 3292
rect 962 3273 969 3277
rect 1001 3272 1008 3280
rect 1615 3237 1624 3249
rect 1686 3253 1692 3258
rect 705 3219 709 3224
rect 1268 3219 1273 3224
<< metal3 >>
rect 344 3317 350 3321
rect 981 3317 1842 3320
rect 981 3313 993 3317
rect 981 3311 988 3313
rect 1839 3292 1842 3317
rect 825 3286 961 3289
rect 825 3283 866 3286
rect 1007 3289 1033 3290
rect 1007 3286 1589 3289
rect 185 3275 188 3279
rect 838 3273 962 3276
rect 1008 3273 1563 3276
rect 40 3236 44 3241
rect 1560 3240 1563 3273
rect 1586 3269 1589 3286
rect 1668 3269 1672 3270
rect 1586 3266 1672 3269
rect 1560 3237 1615 3240
rect 1472 3230 1527 3235
rect 1472 3224 1475 3230
rect 690 3219 705 3224
rect 1273 3219 1475 3224
rect 1524 3222 1527 3230
rect 1533 3222 1537 3228
rect 1524 3219 1537 3222
rect 1525 3218 1537 3219
<< metal4 >>
rect 163 3301 171 3307
rect 810 3298 1648 3302
rect 1644 3283 1648 3298
rect 1644 3279 1659 3283
<< metal5 >>
rect 1465 3239 1546 3244
rect 115 3204 122 3209
rect 1465 3171 1470 3239
rect 1541 3228 1546 3239
rect 1541 3223 1572 3228
rect 1567 3185 1572 3223
rect 859 3166 1470 3171
rect 2766 1630 2932 1634
rect 2766 1606 2770 1630
rect 2928 1626 2932 1630
rect 2766 1598 2774 1606
<< metal6 >>
rect 2920 1541 2925 1553
rect 2920 1536 2930 1541
rect 2925 1317 2930 1536
rect 2824 1312 2930 1317
rect 733 -10 1489 -4
rect 1483 -19 1489 -10
rect 1483 -25 1648 -19
use 7BitDac  7BitDac_0
timestamp 1599268620
transform 1 0 0 0 1 14
box 0 -24 1432 3304
use switchNew  switchNew_0
timestamp 1599222484
transform 1 0 2829 0 1 1550
box 69 -1 187 81
use 7BitDac  7BitDac_1
timestamp 1599268620
transform 1 0 1493 0 1 -5
box 0 -24 1432 3304
<< labels >>
rlabel metal1 16 3249 21 3249 1 R_in8
rlabel metal1 3020 1589 3020 1592 7 V_out8
rlabel metal2 2891 3332 2894 3332 5 D7!
rlabel metal2 2797 3311 2801 3311 1 D6!
rlabel metal3 1586 3289 1589 3289 1 D1!
rlabel metal3 838 3276 841 3276 1 D2!
rlabel space 2623 3240 2626 3240 1 D5!
rlabel metal3 981 3320 988 3320 1 D4!
rlabel metal4 1644 3302 1648 3302 1 D3!
rlabel metal3 40 3241 44 3241 1 D0
rlabel metal3 185 3279 188 3279 1 D2
rlabel metal4 163 3307 171 3307 1 D3
rlabel metal3 344 3321 350 3321 1 D4
rlabel metal2 481 3262 484 3262 1 D5
rlabel metal2 1304 3251 1309 3251 1 D6
rlabel metal3 1533 3228 1537 3228 1 D0!
rlabel metal5 115 3204 122 3204 1 VA
rlabel metal1 2162 -20 2166 -20 1 R_out8
<< end >>
