* SPICE3 file created from 10BitDac.ext - technology: scmos

.model polyResistor R ( TC1=0 TC2=0 RSH=7.7 DEFW=1.E-7 NARROW=0.0 TNOM=27)

.model pfet PMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=4.1589E17 VTH0=-0.3938813 K1=0.5479015 K2=0.0360586 K3=0.0993095 K3B=5.7086622 W0=1E-6 NLX=1.313191E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=0.4911363 DVT1=0.2227356 DVT2=0.1 U0=115.6852975 UA=1.505832E-9 UB=1E-21 UC=-1E-10 VSAT=1.329694E5 A0=1.7590478 AGS=0.3641621 B0=3.427126E-7 B1=1.062928E-6 KETA=0.0134667 A1=0.6859506 A2=0.3506788 RDSW=168.5705677 PRWG=0.5 PRWB=-0.4987371 WR=1 WINT=0 LINT=3.028832E-8 XL=0 XW=-1E-8 DWG=-2.349633E-8 DWB=-7.152486E-9 VOFF=-0.0994037 NFACTOR=1.9424315 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=0.0608072 ETAB=-0.0426148 DSUB=0.7343015 PCLM=3.2579974 PDIBLC1=7.229527E-6 PDIBLC2=0.025389 PDIBLCB=-1E-3 DROUT=0 PSCBE1=1.454878E10 PSCBE2=4.202027E-9 PVAG=15 DELTA=0.01 RSH=7.8 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=6.32E-10 CGSO=6.32E-10 CGBO=1E-12 CJ=1.172138E-3 PB=0.8421173 MJ=0.4109788 CJSW=2.242609E-10 PBSW=0.8 MJSW=0.3752089 CJSWG=4.22E-10 PBSWG=0.8 MJSWG=0.3752089 CF=0 PVTH0=1.888482E-3 PRDSW=11.5315407 PK2=1.559399E-3 WKETA=0.0319301 LKETA=2.955547E-3 PU0=-1.1105313 PUA=-4.62102E-11 PUB=1E-21 PVSAT=50 PETA0=1E-4 PKETA=-4.346368E-3)

.model nfet NMOS (LEVEL=8 VERSION=3.2 TNOM=27 TOX=4.1E-9 XJ=1E-7 NCH=2.3549E17 VTH0=0.3823463 K1=0.5810697 K2=4.774618E-3 K3=0.0431669 K3B=1.1498346 W0=1E-7 NLX=1.910552E-7 DVT0W=0 DVT1W=0 DVT2W=0 DVT0=1.2894824 DVT1=0.3622063 DVT2=0.0713729 U0=280.633249 UA=-1.208537E-9 UB=2.158625E-18 UC=5.342807E-11 VSAT=9.366802E4 A0=1.7593146 AGS=0.3939741 B0=-6.413949E-9 B1=-1E-7 KETA=-5.180424E-4 A1=0 A2=1 RDSW=105.5517558 PRWG=0.5 PRWB=-0.1998871 WR=1 WINT=7.904732E-10 LINT=1.571424E-8 XL=0 XW=-1E-8 DWG=1.297221E-9 DWB=1.479041E-9 VOFF=-0.0955434 NFACTOR=2.4358891 CIT=0 CDSC=2.4E-4 CDSCD=0 CDSCB=0 ETA0=3.104851E-3 ETAB=-2.512384E-5 DSUB=0.0167075 PCLM=0.8073191 PDIBLC1=0.1666161 PDIBLC2=3.112892E-3 PDIBLCB=-0.1 DROUT=0.7875618 PSCBE1=8E10 PSCBE2=9.213635E-10 PVAG=3.85243E-3 DELTA=0.01 RSH=6.7 MOBMOD=1 PRT=0 UTE=-1.5 KT1=-0.11 KT1L=0 KT2=0.022 UA1=4.31E-9 UB1=-7.61E-18 UC1=-5.6E-11 AT=3.3E4 WL=0 WLN=1 WW=0 WWN=1 WWL=0 LL=0 LLN=1 LW=0 LWN=1 LWL=0 CAPMOD=2 XPART=0.5 CGDO=7.08E-10 CGSO=7.08E-10 CGBO=1E-12 CJ=9.68858E-4 PB=0.8 MJ=0.3864502 CJSW=2.512138E-10 PBSW=0.809286 MJSW=0.1060414 CJSWG=3.3E-10 PBSWG=0.809286 MJSWG=0.1060414 CF=0 PVTH0=-1.192722E-3 PRDSW=-5 PK2=6.450505E-5 WKETA=-4.27294E-4 LKETA=-0.0104078 PU0=6.3268729 PUA=2.226552E-11 PUB=0 PVSAT=969.1480157 PETA0=1E-4 PKETA=-1.049509E-3)
.option scale=0.1u

C0 gnd V_out10 3283700.000000fF
M1000 switchNew_0/a_86_24# D9 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=143220 ps=69564
M1001 switchNew_0/a_105_21# switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1002 V_out10 switchNew_0/a_86_24# 9BitDac_0/V_out9 9BitDac_0/V_out9 pfet w=10 l=2
+  ad=140 pd=68 as=210 ps=102
M1003 9BitDac_0/V_out9 switchNew_0/a_105_21# V_out10 gnd nfet w=5 l=2
+  ad=137 pd=104 as=86 ps=64
M1004 switchNew_0/a_86_24# D9 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=71610 ps=49104
M1005 switchNew_0/a_105_21# switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1006 V_out10 switchNew_0/a_86_24# 9BitDac_1/V_out9 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1007 V_out10 switchNew_0/a_105_21# 9BitDac_1/V_out9 V_out10 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1008 9BitDac_1/8BitDac_1/7BitDac_1/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1009 9BitDac_1/8BitDac_1/7BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1010 9BitDac_1/8BitDac_1/7BitDac_1/V_out7 9BitDac_1/8BitDac_1/7BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1011 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 9BitDac_1/8BitDac_1/7BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/V_out7 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1012 9BitDac_1/8BitDac_1/7BitDac_1/switchNew_0/a_86_24# D6 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1013 9BitDac_1/8BitDac_1/7BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1014 9BitDac_1/8BitDac_1/7BitDac_1/V_out7 9BitDac_1/8BitDac_1/7BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1015 9BitDac_1/8BitDac_1/7BitDac_1/V_out7 9BitDac_1/8BitDac_1/7BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 9BitDac_1/8BitDac_1/7BitDac_1/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1016 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1017 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1018 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1019 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1020 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1021 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1022 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1023 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1024 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1025 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1026 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1027 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1028 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1029 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1030 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1031 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1032 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1033 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1034 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1035 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1036 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1037 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1038 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1039 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1040 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1041 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1042 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1043 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1044 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1045 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1046 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1047 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# gnd 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R0 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma gnd polyResistor w=2 l=62
M1048 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1049 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1050 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1051 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1052 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1053 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1054 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1055 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1056 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1057 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1058 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1059 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1060 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1061 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1062 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1065 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1066 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1067 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1068 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1069 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1070 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1071 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1072 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1073 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1074 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1075 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1076 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1077 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1078 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1079 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1080 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1081 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1082 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1083 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1084 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1085 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1086 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1087 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R6 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R7 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1088 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1089 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1090 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1091 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1092 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1093 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1094 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1097 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1098 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1099 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1100 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1101 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1102 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1103 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1104 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1105 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1106 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1107 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1108 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1109 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1110 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1111 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R8 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M1112 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1113 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1114 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1115 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1116 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1117 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1118 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1119 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R9 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R10 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R11 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1120 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1121 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1122 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1123 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1124 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1125 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1126 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1127 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1129 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1130 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1131 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1132 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1133 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1134 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1135 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1136 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1137 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1138 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1139 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1140 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1141 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1142 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1143 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R12 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1144 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1145 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1146 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1147 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1148 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1149 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1150 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1151 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R13 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R14 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R15 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1152 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1153 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1154 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1155 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1156 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1157 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1158 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1159 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1160 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1161 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1162 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1163 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1164 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1165 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1166 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1167 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R16 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M1168 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1169 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1170 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1171 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1172 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1173 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1174 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1175 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R17 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R18 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R19 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1176 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1177 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1178 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1179 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1180 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1181 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1182 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1184 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1185 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1186 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1187 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1188 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1189 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1190 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1191 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1192 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1193 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1194 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1195 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1196 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1197 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1198 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1199 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R20 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1200 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1201 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1202 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1203 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1204 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1205 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1206 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1207 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R21 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R22 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R23 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1208 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1209 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1210 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1211 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1212 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1213 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1214 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1217 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1218 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1219 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1220 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1221 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1222 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1223 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1224 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1225 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1226 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1227 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1228 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1229 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1230 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1231 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R24 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M1232 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1233 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1234 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1235 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1236 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1237 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1238 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1239 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R25 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R26 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R27 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1240 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1241 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1242 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1243 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1244 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1245 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1246 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1247 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1248 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1249 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1250 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1251 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1252 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1253 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1254 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1255 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1256 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1257 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1258 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1259 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1260 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1261 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1262 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1263 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R28 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1264 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1265 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1266 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1267 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1268 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1269 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1270 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1271 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R29 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R30 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R31 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1272 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1273 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1274 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1275 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1276 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1277 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1278 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1279 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1280 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1281 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1282 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1283 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1284 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1285 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1286 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1287 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1288 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1289 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1290 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1291 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1292 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1293 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1294 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1295 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R32 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M1296 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1297 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1298 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1299 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1300 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1301 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1302 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1303 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R33 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R34 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R35 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1304 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1305 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1306 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1307 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1308 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1309 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1310 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1311 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1312 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1313 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1314 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1315 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1316 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1317 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1318 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1319 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1320 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1321 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1322 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1323 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1324 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1325 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1326 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1327 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R36 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1328 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1329 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1330 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1331 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1332 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1333 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1334 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1335 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R37 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R38 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R39 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1336 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1337 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1338 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1339 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1340 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1341 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1342 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1343 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1344 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1345 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1346 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1347 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1348 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1349 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1350 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1351 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1352 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1353 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1354 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1355 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1356 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1357 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1358 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1359 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R40 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M1360 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1361 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1362 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1363 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1364 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1365 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1366 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1367 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R41 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R42 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R43 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1368 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1369 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1370 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1371 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1372 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1373 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1374 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1375 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1376 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1377 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1378 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1379 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1380 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1381 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1382 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1383 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1384 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1385 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1386 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1387 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1388 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1389 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1390 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1391 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R44 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1392 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1393 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1394 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1395 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1396 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1397 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1398 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1399 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R45 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R46 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R47 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1400 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1401 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1402 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1403 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1404 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1405 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1406 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1407 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1408 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1409 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1410 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1411 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1412 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1413 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1414 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1415 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R48 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M1416 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1417 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1418 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1419 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1420 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1421 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1422 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1423 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R49 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R50 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R51 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1424 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1425 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1426 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1427 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1428 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1429 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1430 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1431 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1432 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1433 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1434 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1435 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1436 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1437 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1438 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1439 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1440 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1441 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1442 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1443 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1444 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1445 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1446 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1447 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R52 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1448 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1449 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1450 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1451 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1452 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1453 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1454 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1455 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R53 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R54 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R55 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1456 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1457 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1458 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1459 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1460 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1461 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1462 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1463 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1464 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1465 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1466 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1467 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1468 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1469 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1470 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1471 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1472 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1473 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1474 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1475 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1476 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1477 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1478 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1479 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R56 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M1480 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1481 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1482 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1483 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1484 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1485 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1486 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1487 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R57 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R58 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R59 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1488 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1489 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1490 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1491 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1492 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1493 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1494 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1495 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1496 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1497 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1498 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1499 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1500 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1501 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1502 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1503 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1504 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1505 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1506 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1507 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1508 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1509 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1510 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1511 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R60 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1512 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1513 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1514 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1515 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1516 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1517 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1518 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1519 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R61 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R62 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R63 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/R_in6 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1520 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1521 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1522 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1523 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1524 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1525 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1526 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1527 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1528 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1529 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1530 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1531 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1532 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1533 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1534 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1535 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1536 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1537 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1538 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1539 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1540 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1541 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1542 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1543 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1544 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1545 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1546 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1547 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1548 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1549 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1550 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/R_in6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1551 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/R_in6 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R64 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/R_in6 polyResistor w=2 l=62
M1552 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1553 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1554 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1555 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1556 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1557 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1558 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1559 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R65 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R66 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R67 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1560 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1561 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1562 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1563 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1564 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1565 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1566 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1567 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1568 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1569 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1570 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1571 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1572 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1573 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1574 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1575 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1576 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1577 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1578 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1579 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1580 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1581 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1582 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1583 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R68 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1584 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1585 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1586 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1587 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1588 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1589 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1590 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1591 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R69 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R70 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R71 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1592 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1593 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1594 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1595 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1596 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1597 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1598 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1599 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1600 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1601 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1602 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1603 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1604 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1605 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1606 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1607 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1608 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1609 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1610 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1611 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1612 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1613 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1614 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1615 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R72 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M1616 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1617 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1618 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1619 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1620 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1621 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1622 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1623 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R73 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R74 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R75 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1624 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1625 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1626 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1627 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1628 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1629 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1630 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1631 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1632 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1633 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1634 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1635 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1636 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1637 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1638 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1639 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1640 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1641 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1642 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1643 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1644 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1645 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1646 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1647 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R76 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1648 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1649 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1650 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1651 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1652 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1653 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1654 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1655 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R77 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R78 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R79 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1656 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1657 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1658 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1659 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1660 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1661 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1662 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1663 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1664 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1665 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1666 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1667 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1668 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1669 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1670 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1671 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R80 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M1672 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1673 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1674 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1675 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1676 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1677 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1678 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1679 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R81 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R82 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R83 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1680 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1681 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1682 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1683 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1684 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1685 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1686 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1687 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1688 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1689 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1690 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1691 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1692 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1693 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1694 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1695 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1696 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1697 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1698 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1699 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1700 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1701 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1702 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1703 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R84 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1704 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1705 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1706 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1707 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1708 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1709 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1710 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1711 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R85 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R86 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R87 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1712 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1713 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1714 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1715 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1716 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1717 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1718 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1719 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1720 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1721 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1722 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1723 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1724 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1725 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1726 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1727 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1728 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1729 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1730 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1731 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1732 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1733 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1734 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1735 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R88 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M1736 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1737 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1738 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1739 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1740 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1741 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1742 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1743 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R89 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R90 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R91 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1744 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1745 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1746 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1747 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1748 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1749 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1750 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1751 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1752 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1753 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1754 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1755 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1756 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1757 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1758 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1759 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1760 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1761 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1762 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1763 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1764 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1765 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1766 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1767 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R92 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1768 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1769 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1770 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1771 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1772 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1773 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1774 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1775 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R93 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R94 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R95 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1776 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1777 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1778 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1779 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1780 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1781 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1782 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1783 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1784 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1785 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1786 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1787 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1788 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1789 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1790 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1791 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1792 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1793 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1794 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1795 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1796 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1797 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1798 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1799 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R96 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M1800 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1801 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1802 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1803 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1804 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1805 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1806 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1807 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R97 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R98 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R99 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1808 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1809 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1810 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1811 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1812 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1813 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1814 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1815 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1816 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1817 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1818 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1819 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1820 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1821 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1822 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1823 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1824 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1825 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1826 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1827 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1828 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1829 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1830 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1831 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R100 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1832 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1833 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1834 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1835 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1836 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1837 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1838 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1839 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R101 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R102 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R103 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1840 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1841 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1842 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1843 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1844 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1845 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1846 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1847 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1848 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1849 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1850 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1851 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1852 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1853 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1854 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1855 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1856 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1857 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1858 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1859 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1860 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1861 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1862 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1863 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R104 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M1864 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1865 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1866 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1867 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1868 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1869 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1870 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1871 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R105 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R106 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R107 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1872 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1873 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1874 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1875 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1876 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1877 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1878 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1879 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1880 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1881 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1882 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1883 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1884 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1885 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1886 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1887 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1888 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1889 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1890 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1891 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1892 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1893 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1894 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1895 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R108 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M1896 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1897 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1898 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1899 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1900 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1901 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1902 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1903 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R109 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R110 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R111 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M1904 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1905 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1906 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1907 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1908 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1909 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1910 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1911 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1912 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1913 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1914 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1915 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1916 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1917 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1918 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1919 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R112 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M1920 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1921 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1922 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1923 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1924 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1925 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1926 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1927 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R113 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R114 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R115 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M1928 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1929 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1930 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1931 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1932 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1933 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1934 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1935 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1936 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1937 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1938 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1939 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1940 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1941 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1942 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1943 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1944 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1945 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1946 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1947 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1948 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1949 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1950 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1951 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R116 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M1952 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1953 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1954 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1955 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1956 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1957 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1958 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1959 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R117 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R118 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R119 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M1960 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1961 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1962 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1963 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1964 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1965 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1966 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1967 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1968 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1969 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1970 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M1971 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M1972 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1973 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1974 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M1975 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1976 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1977 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1978 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1979 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1980 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1981 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1982 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1983 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R120 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M1984 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1985 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1986 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M1987 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M1988 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1989 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1990 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M1991 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R121 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R122 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R123 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M1992 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1993 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1994 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M1995 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M1996 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1997 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1998 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M1999 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2000 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2001 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2002 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2003 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2004 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2005 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2006 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2007 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2008 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2009 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2010 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2011 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2012 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2013 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2014 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2015 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R124 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2016 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2017 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2018 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2019 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2020 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2021 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2022 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2023 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R125 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R126 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R127 9BitDac_1/8BitDac_1/7BitDac_1/R_in7 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2024 9BitDac_1/8BitDac_1/switchNew_0/a_86_24# D7 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2025 9BitDac_1/8BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2026 9BitDac_1/8BitDac_1/V_out8 9BitDac_1/8BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/V_out7 9BitDac_1/8BitDac_1/7BitDac_0/V_out7 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2027 9BitDac_1/8BitDac_1/7BitDac_0/V_out7 9BitDac_1/8BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/V_out8 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2028 9BitDac_1/8BitDac_1/switchNew_0/a_86_24# D7 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2029 9BitDac_1/8BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2030 9BitDac_1/8BitDac_1/V_out8 9BitDac_1/8BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/V_out7 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2031 9BitDac_1/8BitDac_1/V_out8 9BitDac_1/8BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/V_out7 9BitDac_1/8BitDac_1/V_out8 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2032 9BitDac_1/8BitDac_1/7BitDac_0/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2033 9BitDac_1/8BitDac_1/7BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2034 9BitDac_1/8BitDac_1/7BitDac_0/V_out7 9BitDac_1/8BitDac_1/7BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2035 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 9BitDac_1/8BitDac_1/7BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/V_out7 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2036 9BitDac_1/8BitDac_1/7BitDac_0/switchNew_0/a_86_24# D6 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2037 9BitDac_1/8BitDac_1/7BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2038 9BitDac_1/8BitDac_1/7BitDac_0/V_out7 9BitDac_1/8BitDac_1/7BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2039 9BitDac_1/8BitDac_1/7BitDac_0/V_out7 9BitDac_1/8BitDac_1/7BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 9BitDac_1/8BitDac_1/7BitDac_0/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2040 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2041 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2042 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2043 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2044 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2045 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2046 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2047 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2048 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2049 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2050 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2051 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2052 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2053 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2054 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2055 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2056 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2057 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2058 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2059 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2060 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2061 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2062 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2063 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2064 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2065 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2066 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2067 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2068 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2069 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2070 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_1/R_in7 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2071 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_1/R_in7 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R128 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_1/R_in7 polyResistor w=2 l=62
M2072 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2073 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2074 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2075 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2076 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2077 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2078 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2079 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R129 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R130 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R131 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2080 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2081 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2082 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2083 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2084 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2085 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2086 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2087 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2088 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2089 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2090 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2091 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2092 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2093 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2094 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2095 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2096 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2097 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2098 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2099 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2100 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2101 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2102 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2103 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R132 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2104 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2105 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2106 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2107 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2108 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2109 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2110 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2111 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R133 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R134 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R135 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2112 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2113 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2114 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2115 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2116 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2117 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2118 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2119 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2120 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2121 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2122 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2123 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2124 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2125 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2126 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2127 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2128 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2129 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2130 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2131 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2132 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2133 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2134 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2135 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R136 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M2136 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2137 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2138 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2139 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2140 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2141 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2142 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2143 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R137 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R138 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R139 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2144 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2145 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2146 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2147 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2148 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2149 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2150 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2151 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2152 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2153 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2154 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2155 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2156 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2157 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2158 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2159 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2160 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2161 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2162 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2163 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2164 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2165 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2166 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2167 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R140 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2168 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2169 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2170 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2171 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2172 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2173 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2174 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2175 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R141 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R142 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R143 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2176 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2177 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2178 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2179 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2180 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2181 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2182 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2183 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2184 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2185 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2186 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2187 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2188 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2189 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2190 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2191 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R144 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M2192 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2193 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2194 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2195 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2196 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2197 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2198 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2199 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R145 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R146 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R147 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2200 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2201 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2202 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2203 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2204 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2205 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2206 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2207 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2208 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2209 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2210 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2211 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2212 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2213 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2214 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2215 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2216 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2217 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2218 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2219 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2220 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2221 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2222 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2223 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R148 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2224 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2225 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2226 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2227 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2228 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2229 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2230 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2231 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R149 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R150 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R151 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2232 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2233 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2234 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2235 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2236 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2237 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2238 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2239 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2240 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2241 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2242 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2243 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2244 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2245 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2246 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2247 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2248 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2249 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2250 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2251 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2252 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2253 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2254 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2255 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R152 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M2256 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2257 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2258 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2259 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2260 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2261 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2262 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2263 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R153 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R154 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R155 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2264 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2265 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2266 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2267 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2268 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2269 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2270 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2271 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2272 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2273 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2274 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2275 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2276 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2277 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2278 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2279 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2280 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2281 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2282 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2283 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2284 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2285 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2286 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2287 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R156 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2288 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2289 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2290 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2291 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2292 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2293 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2294 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2295 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R157 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R158 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R159 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2296 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2297 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2298 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2299 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2300 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2301 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2302 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2303 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2304 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2305 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2306 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2307 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2308 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2309 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2310 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2311 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2312 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2313 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2314 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2315 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2316 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2317 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2318 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2319 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R160 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M2320 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2321 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2322 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2323 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2324 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2325 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2326 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2327 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R161 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R162 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R163 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2328 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2329 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2330 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2331 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2332 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2333 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2334 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2335 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2336 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2337 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2338 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2339 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2340 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2341 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2342 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2343 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2344 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2345 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2346 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2347 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2348 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2349 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2350 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2351 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R164 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2352 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2353 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2354 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2355 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2356 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2357 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2358 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2359 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R165 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R166 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R167 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2360 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2361 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2362 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2363 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2364 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2365 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2366 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2367 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2368 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2369 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2370 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2371 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2372 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2373 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2374 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2375 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2376 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2377 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2378 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2379 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2380 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2381 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2382 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2383 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R168 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M2384 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2385 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2386 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2387 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2388 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2389 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2390 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2391 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R169 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R170 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R171 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2392 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2393 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2394 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2395 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2396 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2397 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2398 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2399 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2400 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2401 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2402 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2403 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2404 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2405 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2406 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2407 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2408 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2409 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2410 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2411 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2412 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2413 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2414 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2415 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R172 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2416 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2417 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2418 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2419 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2420 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2421 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2422 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2423 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R173 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R174 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R175 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2424 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2425 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2426 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2427 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2428 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2429 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2430 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2431 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2432 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2433 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2434 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2435 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2436 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2437 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2438 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2439 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R176 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M2440 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2441 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2442 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2443 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2444 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2445 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2446 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2447 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R177 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R178 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R179 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2448 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2449 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2450 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2451 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2452 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2453 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2454 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2455 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2456 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2457 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2458 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2459 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2460 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2461 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2462 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2463 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2464 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2465 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2466 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2467 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2468 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2469 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2470 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2471 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R180 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2472 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2473 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2474 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2475 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2476 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2477 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2478 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2479 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R181 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R182 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R183 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2480 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2481 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2482 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2483 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2484 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2485 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2486 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2487 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2488 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2489 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2490 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2491 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2492 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2493 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2494 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2495 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2496 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2497 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2498 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2499 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2500 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2501 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2502 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2503 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R184 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M2504 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2505 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2506 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2507 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2508 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2509 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2510 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2511 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R185 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R186 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R187 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2512 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2513 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2514 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2515 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2516 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2517 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2518 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2519 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2520 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2521 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2522 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2523 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2524 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2525 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2526 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2527 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2528 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2529 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2530 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2531 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2532 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2533 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2534 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2535 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R188 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2536 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2537 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2538 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2539 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2540 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2541 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2542 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2543 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R189 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R190 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R191 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/R_in6 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2544 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2545 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2546 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2547 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2548 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2549 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2550 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2551 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2552 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2553 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2554 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2555 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2556 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2557 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2558 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2559 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2560 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2561 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2562 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2563 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2564 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2565 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2566 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2567 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2568 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2569 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2570 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2571 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2572 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2573 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2574 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/R_in6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2575 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/R_in6 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R192 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/R_in6 polyResistor w=2 l=62
M2576 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2577 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2578 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2579 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2580 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2581 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2582 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2583 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R193 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R194 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R195 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2584 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2585 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2586 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2587 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2588 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2589 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2590 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2591 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2592 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2593 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2594 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2595 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2596 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2597 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2598 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2599 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2600 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2601 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2602 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2603 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2604 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2605 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2606 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2607 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R196 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2608 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2609 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2610 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2611 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2612 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2613 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2614 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2615 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R197 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R198 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R199 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2616 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2617 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2618 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2619 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2620 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2621 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2622 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2623 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2624 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2625 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2626 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2627 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2628 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2629 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2630 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2631 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2632 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2633 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2634 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2635 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2636 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2637 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2638 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2639 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R200 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M2640 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2641 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2642 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2643 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2644 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2645 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2646 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2647 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R201 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R202 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R203 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2648 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2649 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2650 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2651 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2652 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2653 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2654 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2655 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2656 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2657 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2658 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2659 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2660 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2661 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2662 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2663 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2664 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2665 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2666 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2667 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2668 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2669 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2670 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2671 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R204 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2672 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2673 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2674 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2675 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2676 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2677 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2678 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2679 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R205 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R206 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R207 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2680 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2681 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2682 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2683 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2684 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2685 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2686 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2687 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2688 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2689 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2690 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2691 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2692 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2693 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2694 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2695 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R208 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M2696 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2697 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2698 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2699 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2700 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2701 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2702 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2703 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R209 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R210 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R211 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2704 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2705 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2706 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2707 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2708 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2709 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2710 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2711 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2712 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2713 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2714 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2715 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2716 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2717 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2718 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2719 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2720 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2721 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2722 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2723 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2724 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2725 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2726 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2727 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R212 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2728 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2729 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2730 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2731 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2732 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2733 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2734 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2735 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R213 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R214 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R215 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2736 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2737 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2738 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2739 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2740 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2741 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2742 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2743 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2744 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2745 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2746 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2747 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2748 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2749 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2750 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2751 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2752 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2753 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2754 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2755 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2756 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2757 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2758 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2759 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R216 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M2760 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2761 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2762 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2763 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2764 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2765 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2766 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2767 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R217 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R218 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R219 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2768 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2769 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2770 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2771 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2772 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2773 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2774 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2775 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2776 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2777 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2778 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2779 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2780 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2781 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2782 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2783 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2784 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2785 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2786 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2787 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2788 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2789 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2790 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2791 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R220 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2792 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2793 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2794 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2795 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2796 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2797 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2798 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2799 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R221 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R222 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R223 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2800 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2801 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2802 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2803 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2804 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2805 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2806 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2807 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2808 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2809 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2810 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2811 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2812 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2813 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2814 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2815 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2816 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2817 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2818 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2819 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2820 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2821 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2822 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2823 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R224 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M2824 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2825 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2826 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2827 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2828 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2829 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2830 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2831 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R225 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R226 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R227 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2832 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2833 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2834 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2835 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2836 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2837 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2838 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2839 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2840 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2841 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2842 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2843 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2844 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2845 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2846 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2847 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2848 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2849 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2850 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2851 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2852 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2853 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2854 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2855 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R228 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2856 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2857 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2858 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2859 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2860 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2861 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2862 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2863 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R229 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R230 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R231 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2864 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2865 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2866 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2867 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2868 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2869 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2870 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2871 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2872 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2873 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2874 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2875 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2876 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2877 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2878 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2879 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2880 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2881 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2882 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2883 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2884 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2885 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2886 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2887 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R232 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M2888 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2889 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2890 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2891 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2892 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2893 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2894 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2895 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R233 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R234 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R235 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M2896 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2897 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2898 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2899 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2900 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2901 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2902 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2903 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2904 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2905 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2906 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2907 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2908 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2909 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2910 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2911 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2912 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2913 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2914 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2915 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2916 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2917 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2918 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2919 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R236 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M2920 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2921 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2922 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2923 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2924 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2925 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2926 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2927 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R237 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R238 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R239 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M2928 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2929 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2930 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2931 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2932 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2933 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2934 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2935 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2936 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2937 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2938 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2939 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2940 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2941 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2942 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2943 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R240 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M2944 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2945 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2946 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2947 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2948 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2949 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2950 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2951 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R241 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R242 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R243 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M2952 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2953 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2954 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2955 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2956 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2957 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2958 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2959 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2960 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2961 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2962 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2963 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2964 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2965 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2966 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2967 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2968 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2969 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2970 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2971 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2972 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2973 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2974 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2975 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R244 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M2976 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2977 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2978 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M2979 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M2980 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2981 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2982 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M2983 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R245 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R246 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R247 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M2984 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2985 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2986 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M2987 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M2988 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2989 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2990 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M2991 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2992 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2993 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M2994 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M2995 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M2996 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2997 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M2998 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M2999 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3000 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3001 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3002 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3003 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3004 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3005 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3006 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3007 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R248 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M3008 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3009 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3010 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3011 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3012 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3013 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3014 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3015 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R249 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R250 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R251 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3016 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3017 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3018 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3019 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3020 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3021 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3022 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3023 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3024 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3025 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3026 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3027 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3028 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3029 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3030 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3031 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3032 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3033 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3034 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3035 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3036 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3037 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3038 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3039 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R252 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3040 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3041 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3042 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3043 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3044 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3045 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3046 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3047 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R253 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R254 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R255 9BitDac_1/8BitDac_1/R_in8 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3048 9BitDac_1/switchNew_0/a_86_24# D8 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3049 9BitDac_1/switchNew_0/a_105_21# 9BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3050 9BitDac_1/V_out9 9BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/V_out8 9BitDac_1/8BitDac_0/V_out8 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3051 9BitDac_1/8BitDac_0/V_out8 9BitDac_1/switchNew_0/a_105_21# 9BitDac_1/V_out9 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3052 9BitDac_1/switchNew_0/a_86_24# D8 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3053 9BitDac_1/switchNew_0/a_105_21# 9BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3054 9BitDac_1/V_out9 9BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_1/V_out8 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3055 9BitDac_1/V_out9 9BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_1/V_out8 9BitDac_1/V_out9 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3056 9BitDac_1/8BitDac_0/7BitDac_1/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3057 9BitDac_1/8BitDac_0/7BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3058 9BitDac_1/8BitDac_0/7BitDac_1/V_out7 9BitDac_1/8BitDac_0/7BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3059 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 9BitDac_1/8BitDac_0/7BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/V_out7 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3060 9BitDac_1/8BitDac_0/7BitDac_1/switchNew_0/a_86_24# D6 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3061 9BitDac_1/8BitDac_0/7BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3062 9BitDac_1/8BitDac_0/7BitDac_1/V_out7 9BitDac_1/8BitDac_0/7BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3063 9BitDac_1/8BitDac_0/7BitDac_1/V_out7 9BitDac_1/8BitDac_0/7BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 9BitDac_1/8BitDac_0/7BitDac_1/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3064 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3065 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3066 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3067 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3068 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3069 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3070 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3071 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3072 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3073 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3074 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3075 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3076 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3077 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3078 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3079 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3080 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3081 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3082 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3083 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3084 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3085 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3086 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3087 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3088 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3089 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3090 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3091 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3092 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3093 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3094 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_1/R_in8 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3095 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_1/R_in8 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R256 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_1/R_in8 polyResistor w=2 l=62
M3096 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3097 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3098 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3099 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3100 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3101 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3102 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3103 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R257 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R258 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R259 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3104 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3105 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3106 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3107 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3108 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3109 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3110 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3111 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3112 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3113 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3114 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3115 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3116 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3117 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3118 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3119 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3120 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3121 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3122 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3123 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3124 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3125 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3126 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3127 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R260 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3128 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3129 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3130 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3131 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3132 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3133 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3134 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3135 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R261 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R262 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R263 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3136 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3137 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3138 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3139 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3140 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3141 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3142 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3143 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3144 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3145 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3146 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3147 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3148 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3149 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3150 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3151 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3152 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3153 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3154 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3155 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3156 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3157 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3158 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3159 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R264 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M3160 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3161 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3162 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3163 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3164 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3165 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3166 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3167 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R265 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R266 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R267 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3168 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3169 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3170 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3171 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3172 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3173 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3174 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3175 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3176 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3177 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3178 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3179 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3180 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3181 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3182 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3183 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3184 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3185 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3186 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3187 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3188 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3189 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3190 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3191 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R268 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3192 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3193 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3194 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3195 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3196 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3197 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3198 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3199 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R269 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R270 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R271 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3200 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3201 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3202 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3203 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3204 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3205 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3206 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3207 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3208 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3209 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3210 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3211 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3212 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3213 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3214 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3215 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R272 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M3216 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3217 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3218 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3219 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3220 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3221 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3222 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3223 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R273 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R274 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R275 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3224 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3225 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3226 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3227 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3228 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3229 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3230 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3231 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3232 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3233 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3234 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3235 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3236 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3237 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3238 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3239 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3240 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3241 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3242 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3243 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3244 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3245 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3246 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3247 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R276 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3248 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3249 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3250 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3251 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3252 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3253 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3254 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3255 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R277 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R278 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R279 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3256 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3257 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3258 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3259 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3260 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3261 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3262 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3263 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3264 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3265 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3266 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3267 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3268 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3269 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3270 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3271 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3272 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3273 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3274 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3275 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3276 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3277 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3278 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3279 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R280 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M3280 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3281 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3282 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3283 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3284 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3285 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3286 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3287 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R281 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R282 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R283 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3288 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3289 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3290 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3291 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3292 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3293 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3294 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3295 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3296 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3297 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3298 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3299 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3300 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3301 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3302 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3303 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3304 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3305 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3306 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3307 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3308 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3309 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3310 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3311 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R284 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3312 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3313 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3314 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3315 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3316 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3317 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3318 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3319 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R285 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R286 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R287 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3320 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3321 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3322 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3323 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3324 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3325 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3326 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3327 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3328 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3329 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3330 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3331 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3332 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3333 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3334 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3335 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3336 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3337 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3338 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3339 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3340 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3341 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3342 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3343 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R288 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M3344 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3345 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3346 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3347 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3348 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3349 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3350 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3351 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R289 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R290 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R291 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3352 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3353 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3354 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3355 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3356 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3357 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3358 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3359 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3360 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3361 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3362 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3363 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3364 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3365 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3366 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3367 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3368 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3369 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3370 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3371 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3372 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3373 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3374 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3375 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R292 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3376 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3377 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3378 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3379 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3380 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3381 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3382 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3383 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R293 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R294 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R295 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3384 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3385 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3386 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3387 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3388 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3389 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3390 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3391 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3392 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3393 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3394 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3395 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3396 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3397 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3398 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3399 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3400 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3401 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3402 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3403 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3404 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3405 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3406 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3407 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R296 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M3408 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3409 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3410 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3411 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3412 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3413 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3414 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3415 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R297 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R298 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R299 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3416 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3417 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3418 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3419 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3420 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3421 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3422 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3423 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3424 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3425 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3426 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3427 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3428 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3429 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3430 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3431 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3432 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3433 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3434 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3435 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3436 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3437 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3438 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3439 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R300 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3440 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3441 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3442 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3443 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3444 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3445 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3446 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3447 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R301 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R302 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R303 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3448 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3449 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3450 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3451 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3452 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3453 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3454 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3455 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3456 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3457 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3458 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3459 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3460 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3461 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3462 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3463 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R304 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M3464 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3465 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3466 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3467 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3468 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3469 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3470 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3471 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R305 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R306 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R307 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3472 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3473 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3474 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3475 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3476 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3477 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3478 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3479 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3480 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3481 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3482 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3483 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3484 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3485 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3486 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3487 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3488 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3489 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3490 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3491 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3492 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3493 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3494 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3495 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R308 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3496 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3497 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3498 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3499 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3500 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3501 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3502 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3503 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R309 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R310 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R311 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3504 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3505 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3506 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3507 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3508 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3509 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3510 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3511 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3512 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3513 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3514 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3515 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3516 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3517 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3518 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3519 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3520 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3521 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3522 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3523 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3524 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3525 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3526 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3527 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R312 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M3528 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3529 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3530 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3531 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3532 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3533 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3534 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3535 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R313 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R314 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R315 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3536 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3537 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3538 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3539 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3540 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3541 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3542 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3543 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3544 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3545 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3546 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3547 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3548 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3549 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3550 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3551 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3552 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3553 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3554 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3555 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3556 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3557 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3558 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3559 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R316 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3560 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3561 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3562 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3563 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3564 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3565 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3566 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3567 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R317 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R318 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R319 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/R_in6 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3568 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3569 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3570 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3571 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3572 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3573 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3574 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3575 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3576 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3577 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3578 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3579 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3580 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3581 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3582 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3583 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3584 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3585 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3586 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3587 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3588 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3589 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3590 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3591 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3592 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3593 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3594 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3595 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3596 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3597 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3598 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/R_in6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3599 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/R_in6 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R320 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/R_in6 polyResistor w=2 l=62
M3600 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3601 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3602 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3603 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3604 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3605 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3606 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3607 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R321 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R322 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R323 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3608 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3609 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3610 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3611 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3612 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3613 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3614 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3615 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3616 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3617 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3618 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3619 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3620 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3621 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3622 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3623 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3624 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3625 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3626 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3627 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3628 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3629 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3630 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3631 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R324 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3632 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3633 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3634 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3635 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3636 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3637 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3638 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3639 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R325 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R326 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R327 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3640 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3641 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3642 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3643 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3644 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3645 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3646 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3647 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3648 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3649 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3650 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3651 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3652 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3653 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3654 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3655 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3656 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3657 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3658 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3659 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3660 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3661 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3662 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3663 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R328 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M3664 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3665 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3666 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3667 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3668 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3669 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3670 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3671 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R329 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R330 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R331 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3672 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3673 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3674 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3675 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3676 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3677 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3678 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3679 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3680 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3681 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3682 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3683 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3684 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3685 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3686 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3687 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3688 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3689 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3690 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3691 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3692 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3693 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3694 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3695 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R332 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3696 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3697 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3698 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3699 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3700 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3701 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3702 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3703 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R333 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R334 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R335 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3704 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3705 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3706 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3707 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3708 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3709 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3710 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3711 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3712 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3713 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3714 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3715 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3716 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3717 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3718 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3719 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R336 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M3720 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3721 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3722 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3723 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3724 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3725 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3726 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3727 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R337 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R338 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R339 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3728 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3729 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3730 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3731 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3732 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3733 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3734 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3735 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3736 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3737 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3738 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3739 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3740 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3741 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3742 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3743 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3744 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3745 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3746 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3747 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3748 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3749 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3750 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3751 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R340 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3752 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3753 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3754 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3755 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3756 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3757 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3758 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3759 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R341 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R342 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R343 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3760 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3761 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3762 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3763 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3764 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3765 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3766 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3767 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3768 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3769 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3770 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3771 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3772 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3773 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3774 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3775 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3776 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3777 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3778 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3779 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3780 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3781 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3782 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3783 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R344 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M3784 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3785 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3786 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3787 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3788 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3789 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3790 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3791 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R345 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R346 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R347 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3792 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3793 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3794 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3795 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3796 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3797 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3798 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3799 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3800 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3801 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3802 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3803 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3804 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3805 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3806 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3807 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3808 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3809 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3810 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3811 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3812 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3813 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3814 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3815 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R348 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3816 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3817 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3818 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3819 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3820 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3821 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3822 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3823 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R349 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R350 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R351 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3824 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3825 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3826 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3827 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3828 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3829 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3830 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3831 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3832 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3833 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3834 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3835 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3836 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3837 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3838 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3839 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3840 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3841 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3842 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3843 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3844 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3845 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3846 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3847 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R352 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M3848 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3849 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3850 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3851 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3852 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3853 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3854 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3855 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R353 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R354 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R355 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3856 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3857 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3858 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3859 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3860 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3861 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3862 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3863 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3864 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3865 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3866 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3867 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3868 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3869 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3870 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3871 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3872 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3873 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3874 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3875 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3876 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3877 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3878 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3879 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R356 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M3880 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3881 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3882 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3883 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3884 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3885 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3886 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3887 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R357 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R358 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R359 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M3888 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3889 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3890 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3891 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3892 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3893 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3894 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3895 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3896 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3897 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3898 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3899 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3900 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3901 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3902 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3903 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3904 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3905 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3906 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3907 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3908 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3909 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3910 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3911 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R360 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M3912 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3913 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3914 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3915 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3916 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3917 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3918 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3919 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R361 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R362 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R363 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M3920 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3921 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3922 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3923 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3924 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3925 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3926 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3927 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3928 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3929 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3930 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3931 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3932 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3933 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3934 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3935 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3936 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3937 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3938 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3939 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3940 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3941 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3942 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3943 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R364 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M3944 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3945 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3946 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3947 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3948 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3949 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3950 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3951 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R365 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R366 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R367 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M3952 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3953 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3954 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3955 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3956 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3957 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3958 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3959 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3960 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3961 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3962 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3963 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3964 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3965 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3966 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3967 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R368 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M3968 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3969 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3970 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3971 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3972 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3973 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3974 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3975 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R369 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R370 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R371 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M3976 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3977 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3978 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M3979 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M3980 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3981 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3982 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M3983 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3984 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3985 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3986 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3987 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M3988 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3989 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3990 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M3991 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M3992 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3993 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M3994 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M3995 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M3996 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3997 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M3998 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M3999 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R372 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4000 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4001 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4002 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4003 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4004 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4005 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4006 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4007 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R373 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R374 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R375 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4008 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4009 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4010 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4011 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4012 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4013 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4014 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4015 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4016 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4017 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4018 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4019 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4020 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4021 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4022 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4023 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4024 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4025 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4026 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4027 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4028 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4029 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4030 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4031 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R376 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M4032 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4033 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4034 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4035 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4036 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4037 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4038 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4039 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R377 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R378 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R379 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4040 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4041 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4042 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4043 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4044 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4045 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4046 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4047 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4048 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4049 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4050 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4051 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4052 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4053 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4054 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4055 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4056 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4057 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4058 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4059 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4060 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4061 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4062 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4063 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R380 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4064 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4065 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4066 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4067 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4068 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4069 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4070 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4071 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R381 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R382 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R383 9BitDac_1/8BitDac_0/7BitDac_1/R_in7 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4072 9BitDac_1/8BitDac_0/switchNew_0/a_86_24# D7 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4073 9BitDac_1/8BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4074 9BitDac_1/8BitDac_0/V_out8 9BitDac_1/8BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/V_out7 9BitDac_1/8BitDac_0/7BitDac_0/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4075 9BitDac_1/8BitDac_0/7BitDac_0/V_out7 9BitDac_1/8BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/V_out8 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4076 9BitDac_1/8BitDac_0/switchNew_0/a_86_24# D7 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4077 9BitDac_1/8BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4078 9BitDac_1/8BitDac_0/V_out8 9BitDac_1/8BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/V_out7 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4079 9BitDac_1/8BitDac_0/V_out8 9BitDac_1/8BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/V_out7 9BitDac_1/8BitDac_0/V_out8 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4080 9BitDac_1/8BitDac_0/7BitDac_0/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4081 9BitDac_1/8BitDac_0/7BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4082 9BitDac_1/8BitDac_0/7BitDac_0/V_out7 9BitDac_1/8BitDac_0/7BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4083 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 9BitDac_1/8BitDac_0/7BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/V_out7 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4084 9BitDac_1/8BitDac_0/7BitDac_0/switchNew_0/a_86_24# D6 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4085 9BitDac_1/8BitDac_0/7BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4086 9BitDac_1/8BitDac_0/7BitDac_0/V_out7 9BitDac_1/8BitDac_0/7BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4087 9BitDac_1/8BitDac_0/7BitDac_0/V_out7 9BitDac_1/8BitDac_0/7BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 9BitDac_1/8BitDac_0/7BitDac_0/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4088 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4089 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4090 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4091 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4092 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4093 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4094 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4095 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4096 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4097 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4098 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4099 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4100 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4101 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4102 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4103 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4104 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4105 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4106 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4107 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4108 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4109 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4110 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4111 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4112 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4113 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4114 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4115 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4116 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4117 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4118 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_1/R_in7 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4119 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_1/R_in7 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R384 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_1/R_in7 polyResistor w=2 l=62
M4120 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4121 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4122 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4123 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4124 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4125 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4126 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4127 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R385 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R386 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R387 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4128 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4129 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4130 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4131 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4132 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4133 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4134 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4135 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4136 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4137 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4138 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4139 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4140 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4141 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4142 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4143 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4144 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4145 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4146 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4147 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4148 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4149 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4150 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4151 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R388 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4152 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4153 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4154 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4155 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4156 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4157 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4158 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4159 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R389 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R390 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R391 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4160 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4161 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4162 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4163 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4164 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4165 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4166 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4167 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4168 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4169 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4170 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4171 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4172 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4173 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4174 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4175 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4176 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4177 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4178 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4179 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4180 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4181 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4182 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4183 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R392 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M4184 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4185 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4186 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4187 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4188 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4189 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4190 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4191 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R393 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R394 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R395 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4192 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4193 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4194 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4195 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4196 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4197 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4198 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4199 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4200 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4201 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4202 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4203 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4204 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4205 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4206 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4207 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4208 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4209 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4210 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4211 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4212 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4213 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4214 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4215 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R396 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4216 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4217 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4218 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4219 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4220 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4221 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4222 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4223 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R397 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R398 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R399 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4224 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4225 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4226 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4227 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4228 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4229 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4230 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4231 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4232 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4233 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4234 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4235 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4236 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4237 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4238 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4239 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R400 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M4240 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4241 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4242 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4243 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4244 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4245 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4246 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4247 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R401 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R402 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R403 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4248 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4249 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4250 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4251 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4252 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4253 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4254 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4255 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4256 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4257 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4258 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4259 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4260 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4261 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4262 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4263 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4264 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4265 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4266 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4267 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4268 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4269 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4270 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4271 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R404 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4272 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4273 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4274 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4275 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4276 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4277 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4278 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4279 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R405 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R406 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R407 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4280 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4281 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4282 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4283 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4284 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4285 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4286 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4287 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4288 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4289 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4290 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4291 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4292 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4293 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4294 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4295 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4296 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4297 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4298 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4299 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4300 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4301 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4302 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4303 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R408 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M4304 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4305 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4306 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4307 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4308 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4309 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4310 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4311 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R409 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R410 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R411 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4312 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4313 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4314 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4315 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4316 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4317 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4318 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4319 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4320 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4321 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4322 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4323 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4324 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4325 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4326 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4327 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4328 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4329 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4330 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4331 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4332 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4333 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4334 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4335 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R412 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4336 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4337 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4338 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4339 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4340 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4341 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4342 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4343 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R413 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R414 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R415 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4344 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4345 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4346 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4347 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4348 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4349 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4350 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4351 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4352 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4353 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4354 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4355 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4356 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4357 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4358 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4359 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4360 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4361 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4362 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4363 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4364 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4365 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4366 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4367 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R416 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M4368 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4369 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4370 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4371 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4372 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4373 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4374 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4375 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R417 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R418 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R419 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4376 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4377 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4378 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4379 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4380 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4381 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4382 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4383 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4384 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4385 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4386 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4387 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4388 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4389 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4390 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4391 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4392 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4393 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4394 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4395 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4396 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4397 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4398 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4399 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R420 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4400 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4401 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4402 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4403 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4404 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4405 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4406 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4407 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R421 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R422 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R423 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4408 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4409 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4410 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4411 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4412 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4413 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4414 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4415 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4416 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4417 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4418 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4419 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4420 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4421 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4422 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4423 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4424 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4425 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4426 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4427 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4428 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4429 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4430 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4431 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R424 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M4432 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4433 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4434 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4435 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4436 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4437 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4438 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4439 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R425 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R426 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R427 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4440 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4441 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4442 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4443 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4444 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4445 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4446 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4447 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4448 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4449 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4450 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4451 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4452 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4453 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4454 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4455 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4456 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4457 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4458 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4459 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4460 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4461 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4462 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4463 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R428 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4464 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4465 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4466 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4467 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4468 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4469 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4470 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4471 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R429 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R430 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R431 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4472 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4473 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4474 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4475 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4476 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4477 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4478 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4479 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4480 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4481 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4482 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4483 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4484 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4485 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4486 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4487 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R432 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M4488 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4489 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4490 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4491 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4492 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4493 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4494 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4495 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R433 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R434 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R435 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4496 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4497 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4498 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4499 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4500 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4501 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4502 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4503 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4504 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4505 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4506 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4507 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4508 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4509 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4510 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4511 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4512 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4513 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4514 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4515 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4516 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4517 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4518 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4519 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R436 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4520 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4521 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4522 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4523 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4524 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4525 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4526 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4527 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R437 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R438 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R439 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4528 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4529 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4530 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4531 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4532 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4533 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4534 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4535 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4536 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4537 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4538 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4539 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4540 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4541 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4542 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4543 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4544 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4545 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4546 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4547 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4548 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4549 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4550 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4551 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R440 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M4552 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4553 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4554 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4555 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4556 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4557 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4558 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4559 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R441 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R442 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R443 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4560 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4561 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4562 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4563 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4564 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4565 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4566 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4567 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4568 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4569 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4570 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4571 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4572 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4573 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4574 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4575 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4576 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4577 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4578 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4579 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4580 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4581 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4582 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4583 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R444 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4584 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4585 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4586 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4587 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4588 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4589 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4590 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4591 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R445 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R446 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R447 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/R_in6 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4592 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4593 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4594 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4595 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4596 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4597 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4598 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4599 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4600 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4601 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4602 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4603 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4604 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4605 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4606 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4607 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4608 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4609 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4610 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4611 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4612 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4613 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4614 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4615 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4616 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4617 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4618 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4619 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4620 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4621 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4622 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/R_in6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4623 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/R_in6 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R448 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/R_in6 polyResistor w=2 l=62
M4624 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4625 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4626 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4627 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4628 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4629 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4630 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4631 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R449 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R450 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R451 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4632 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4633 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4634 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4635 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4636 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4637 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4638 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4639 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4640 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4641 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4642 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4643 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4644 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4645 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4646 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4647 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4648 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4649 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4650 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4651 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4652 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4653 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4654 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4655 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R452 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4656 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4657 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4658 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4659 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4660 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4661 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4662 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4663 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R453 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R454 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R455 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4664 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4665 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4666 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4667 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4668 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4669 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4670 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4671 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4672 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4673 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4674 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4675 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4676 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4677 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4678 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4679 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4680 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4681 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4682 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4683 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4684 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4685 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4686 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4687 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R456 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M4688 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4689 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4690 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4691 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4692 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4693 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4694 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4695 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R457 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R458 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R459 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4696 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4697 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4698 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4699 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4700 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4701 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4702 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4703 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4704 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4705 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4706 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4707 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4708 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4709 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4710 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4711 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4712 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4713 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4714 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4715 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4716 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4717 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4718 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4719 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R460 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4720 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4721 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4722 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4723 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4724 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4725 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4726 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4727 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R461 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R462 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R463 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4728 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4729 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4730 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4731 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4732 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4733 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4734 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4735 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4736 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4737 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4738 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4739 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4740 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4741 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4742 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4743 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R464 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M4744 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4745 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4746 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4747 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4748 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4749 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4750 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4751 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R465 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R466 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R467 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4752 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4753 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4754 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4755 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4756 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4757 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4758 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4759 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4760 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4761 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4762 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4763 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4764 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4765 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4766 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4767 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4768 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4769 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4770 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4771 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4772 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4773 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4774 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4775 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R468 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4776 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4777 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4778 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4779 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4780 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4781 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4782 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4783 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R469 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R470 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R471 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4784 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4785 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4786 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4787 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4788 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4789 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4790 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4791 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4792 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4793 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4794 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4795 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4796 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4797 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4798 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4799 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4800 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4801 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4802 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4803 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4804 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4805 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4806 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4807 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R472 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M4808 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4809 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4810 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4811 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4812 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4813 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4814 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4815 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R473 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R474 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R475 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4816 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4817 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4818 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4819 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4820 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4821 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4822 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4823 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4824 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4825 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4826 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4827 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4828 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4829 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4830 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4831 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4832 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4833 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4834 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4835 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4836 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4837 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4838 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4839 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R476 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4840 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4841 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4842 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4843 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4844 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4845 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4846 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4847 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R477 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R478 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R479 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4848 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4849 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4850 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4851 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4852 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4853 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4854 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4855 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4856 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4857 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4858 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4859 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4860 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4861 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4862 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4863 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4864 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4865 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4866 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4867 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4868 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4869 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4870 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4871 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R480 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M4872 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4873 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4874 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4875 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4876 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4877 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4878 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4879 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R481 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R482 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R483 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M4880 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4881 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4882 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4883 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4884 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4885 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4886 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4887 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4888 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4889 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4890 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4891 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4892 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4893 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4894 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4895 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4896 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4897 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4898 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4899 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4900 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4901 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4902 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4903 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R484 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M4904 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4905 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4906 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4907 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4908 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4909 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4910 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4911 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R485 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R486 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R487 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M4912 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4913 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4914 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4915 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4916 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4917 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4918 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4919 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4920 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4921 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4922 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4923 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4924 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4925 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4926 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4927 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4928 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4929 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4930 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4931 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4932 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4933 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4934 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4935 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R488 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M4936 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4937 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4938 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4939 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4940 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4941 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4942 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4943 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R489 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R490 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R491 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M4944 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4945 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4946 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4947 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4948 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4949 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4950 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M4951 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4952 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4953 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4954 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4955 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M4956 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4957 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4958 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4959 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4960 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4961 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4962 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4963 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4964 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4965 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4966 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4967 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R492 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M4968 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4969 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4970 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4971 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4972 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4973 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4974 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4975 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R493 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R494 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R495 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M4976 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4977 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4978 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M4979 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M4980 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4981 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4982 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M4983 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M4984 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4985 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4986 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4987 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4988 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4989 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4990 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4991 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R496 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M4992 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4993 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M4994 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M4995 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M4996 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4997 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M4998 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M4999 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R497 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R498 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R499 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M5000 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5001 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5002 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5003 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5004 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5005 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5006 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5007 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5008 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5009 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5010 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5011 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5012 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5013 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5014 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5015 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5016 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5017 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5018 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5019 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5020 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5021 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5022 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5023 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R500 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M5024 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5025 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5026 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5027 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5028 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5029 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5030 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5031 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R501 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R502 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R503 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M5032 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5033 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5034 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5035 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5036 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5037 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5038 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5039 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5040 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5041 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5042 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5043 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5044 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5045 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5046 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5047 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5048 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5049 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5050 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5051 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5052 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5053 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5054 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5055 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R504 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M5056 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5057 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5058 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5059 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5060 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5061 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5062 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5063 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R505 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R506 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R507 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M5064 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5065 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5066 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5067 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5068 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5069 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5070 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5071 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5072 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5073 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5074 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5075 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5076 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5077 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5078 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5079 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5080 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5081 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5082 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5083 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5084 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5085 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5086 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5087 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R508 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M5088 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5089 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5090 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5091 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5092 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5093 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5094 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5095 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R509 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R510 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R511 9BitDac_1/R_in9 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M5096 9BitDac_0/8BitDac_1/7BitDac_1/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5097 9BitDac_0/8BitDac_1/7BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5098 9BitDac_0/8BitDac_1/7BitDac_1/V_out7 9BitDac_0/8BitDac_1/7BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5099 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 9BitDac_0/8BitDac_1/7BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/V_out7 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5100 9BitDac_0/8BitDac_1/7BitDac_1/switchNew_0/a_86_24# D6 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5101 9BitDac_0/8BitDac_1/7BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5102 9BitDac_0/8BitDac_1/7BitDac_1/V_out7 9BitDac_0/8BitDac_1/7BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5103 9BitDac_0/8BitDac_1/7BitDac_1/V_out7 9BitDac_0/8BitDac_1/7BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 9BitDac_0/8BitDac_1/7BitDac_1/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5104 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5105 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5106 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5107 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5108 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5109 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5110 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5111 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5112 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5113 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5114 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5115 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5116 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5117 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5118 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5119 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5120 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5121 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5122 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5123 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5124 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5125 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5126 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5127 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5128 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5129 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5130 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5131 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5132 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5133 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5134 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_1/R_in9 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5135 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_1/R_in9 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R512 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_1/R_in9 polyResistor w=2 l=62
M5136 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5137 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5138 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5139 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5140 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5141 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5142 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5143 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R513 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R514 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R515 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M5144 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5145 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5146 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5147 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5148 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5149 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5150 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5151 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5152 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5153 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5154 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5155 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5156 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5157 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5158 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5159 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5160 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5161 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5162 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5163 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5164 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5165 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5166 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5167 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R516 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M5168 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5169 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5170 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5171 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5172 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5173 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5174 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5175 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R517 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R518 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R519 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M5176 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5177 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5178 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5179 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5180 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5181 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5182 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5183 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5184 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5185 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5186 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5187 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5188 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5189 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5190 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5191 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5192 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5193 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5194 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5195 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5196 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5197 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5198 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5199 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R520 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M5200 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5201 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5202 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5203 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5204 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5205 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5206 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5207 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R521 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R522 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R523 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M5208 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5209 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5210 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5211 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5212 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5213 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5214 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5215 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5216 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5217 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5218 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5219 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5220 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5221 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5222 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5223 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5224 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5225 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5226 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5227 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5228 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5229 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5230 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5231 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R524 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M5232 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5233 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5234 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5235 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5236 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5237 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5238 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5239 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R525 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R526 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R527 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M5240 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5241 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5242 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5243 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5244 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5245 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5246 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5247 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5248 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5249 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5250 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5251 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5252 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5253 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5254 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5255 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R528 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M5256 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5257 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5258 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5259 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5260 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5261 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5262 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5263 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R529 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R530 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R531 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M5264 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5265 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5266 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5267 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5268 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5269 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5270 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5271 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5272 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5273 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5274 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5275 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5276 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5277 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5278 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5279 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5280 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5281 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5282 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5283 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5284 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5285 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5286 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5287 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R532 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M5288 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5289 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5290 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5291 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5292 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5293 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5294 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5295 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R533 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R534 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R535 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M5296 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5297 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5298 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5299 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5300 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5301 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5302 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5303 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5304 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5305 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5306 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5307 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5308 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5309 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5310 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5311 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5312 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5313 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5314 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5315 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5316 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5317 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5318 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5319 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R536 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M5320 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5321 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5322 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5323 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5324 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5325 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5326 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5327 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R537 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R538 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R539 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M5328 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5329 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5330 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5331 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5332 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5333 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5334 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5335 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5336 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5337 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5338 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5339 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5340 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5341 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5342 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5343 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5344 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5345 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5346 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5347 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5348 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5349 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5350 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5351 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R540 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M5352 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5353 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5354 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5355 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5356 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5357 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5358 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5359 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R541 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R542 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R543 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M5360 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5361 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5362 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5363 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5364 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5365 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5366 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5367 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5368 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5369 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5370 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5371 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5372 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5373 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5374 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5375 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5376 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5377 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5378 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5379 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5380 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5381 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5382 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5383 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R544 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M5384 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5385 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5386 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5387 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5388 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5389 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5390 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5391 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R545 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R546 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R547 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M5392 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5393 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5394 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5395 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5396 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5397 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5398 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5399 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5400 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5401 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5402 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5403 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5404 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5405 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5406 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5407 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5408 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5409 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5410 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5411 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5412 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5413 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5414 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5415 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R548 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M5416 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5417 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5418 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5419 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5420 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5421 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5422 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5423 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R549 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R550 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R551 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M5424 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5425 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5426 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5427 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5428 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5429 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5430 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5431 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5432 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5433 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5434 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5435 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5436 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5437 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5438 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5439 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5440 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5441 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5442 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5443 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5444 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5445 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5446 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5447 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R552 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M5448 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5449 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5450 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5451 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5452 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5453 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5454 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5455 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R553 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R554 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R555 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M5456 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5457 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5458 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5459 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5460 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5461 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5462 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5463 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5464 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5465 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5466 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5467 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5468 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5469 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5470 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5471 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5472 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5473 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5474 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5475 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5476 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5477 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5478 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5479 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R556 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M5480 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5481 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5482 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5483 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5484 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5485 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5486 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5487 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R557 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R558 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R559 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M5488 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5489 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5490 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5491 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5492 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5493 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5494 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5495 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5496 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5497 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5498 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5499 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5500 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5501 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5502 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5503 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R560 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M5504 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5505 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5506 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5507 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5508 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5509 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5510 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5511 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R561 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R562 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R563 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M5512 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5513 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5514 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5515 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5516 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5517 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5518 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5519 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5520 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5521 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5522 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5523 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5524 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5525 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5526 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5527 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5528 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5529 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5530 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5531 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5532 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5533 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5534 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5535 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R564 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M5536 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5537 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5538 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5539 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5540 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5541 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5542 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5543 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R565 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R566 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R567 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M5544 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5545 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5546 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5547 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5548 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5549 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5550 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5551 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5552 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5553 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5554 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5555 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5556 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5557 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5558 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5559 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5560 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5561 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5562 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5563 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5564 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5565 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5566 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5567 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R568 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M5568 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5569 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5570 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5571 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5572 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5573 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5574 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5575 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R569 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R570 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R571 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M5576 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5577 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5578 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5579 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5580 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5581 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5582 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5583 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5584 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5585 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5586 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5587 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5588 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5589 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5590 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5591 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5592 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5593 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5594 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5595 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5596 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5597 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5598 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5599 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R572 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M5600 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5601 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5602 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5603 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5604 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5605 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5606 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5607 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R573 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R574 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R575 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/R_in6 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M5608 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5609 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5610 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5611 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5612 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5613 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5614 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5615 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5616 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5617 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5618 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5619 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5620 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5621 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5622 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5623 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5624 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5625 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5626 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5627 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5628 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5629 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5630 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5631 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5632 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5633 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5634 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5635 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5636 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5637 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5638 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/R_in6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5639 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/R_in6 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R576 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/R_in6 polyResistor w=2 l=62
M5640 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5641 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5642 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5643 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5644 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5645 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5646 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5647 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R577 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R578 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R579 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M5648 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5649 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5650 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5651 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5652 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5653 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5654 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5655 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5656 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5657 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5658 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5659 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5660 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5661 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5662 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5663 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5664 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5665 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5666 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5667 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5668 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5669 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5670 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5671 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R580 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M5672 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5673 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5674 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5675 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5676 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5677 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5678 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5679 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R581 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R582 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R583 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M5680 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5681 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5682 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5683 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5684 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5685 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5686 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5687 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5688 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5689 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5690 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5691 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5692 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5693 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5694 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5695 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5696 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5697 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5698 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5699 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5700 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5701 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5702 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5703 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R584 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M5704 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5705 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5706 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5707 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5708 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5709 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5710 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5711 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R585 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R586 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R587 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M5712 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5713 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5714 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5715 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5716 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5717 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5718 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5719 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5720 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5721 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5722 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5723 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5724 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5725 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5726 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5727 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5728 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5729 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5730 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5731 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5732 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5733 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5734 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5735 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R588 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M5736 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5737 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5738 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5739 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5740 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5741 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5742 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5743 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R589 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R590 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R591 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M5744 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5745 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5746 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5747 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5748 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5749 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5750 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5751 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5752 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5753 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5754 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5755 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5756 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5757 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5758 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5759 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R592 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M5760 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5761 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5762 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5763 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5764 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5765 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5766 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5767 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R593 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R594 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R595 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M5768 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5769 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5770 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5771 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5772 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5773 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5774 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5775 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5776 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5777 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5778 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5779 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5780 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5781 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5782 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5783 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5784 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5785 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5786 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5787 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5788 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5789 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5790 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5791 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R596 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M5792 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5793 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5794 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5795 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5796 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5797 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5798 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5799 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R597 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R598 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R599 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M5800 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5801 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5802 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5803 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5804 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5805 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5806 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5807 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5808 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5809 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5810 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5811 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5812 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5813 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5814 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5815 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5816 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5817 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5818 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5819 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5820 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5821 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5822 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5823 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R600 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M5824 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5825 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5826 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5827 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5828 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5829 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5830 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5831 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R601 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R602 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R603 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M5832 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5833 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5834 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5835 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5836 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5837 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5838 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5839 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5840 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5841 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5842 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5843 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5844 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5845 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5846 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5847 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5848 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5849 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5850 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5851 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5852 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5853 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5854 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5855 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R604 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M5856 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5857 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5858 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5859 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5860 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5861 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5862 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5863 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R605 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R606 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R607 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M5864 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5865 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5866 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5867 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5868 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5869 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5870 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5871 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5872 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5873 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5874 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5875 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5876 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5877 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5878 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5879 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5880 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5881 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5882 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5883 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5884 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5885 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5886 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5887 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R608 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M5888 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5889 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5890 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5891 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5892 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5893 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5894 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5895 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R609 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R610 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R611 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M5896 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5897 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5898 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5899 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5900 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5901 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5902 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5903 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5904 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5905 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5906 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5907 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5908 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5909 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5910 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5911 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5912 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5913 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5914 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5915 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5916 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5917 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5918 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5919 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R612 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M5920 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5921 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5922 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5923 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5924 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5925 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5926 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5927 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R613 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R614 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R615 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M5928 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5929 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5930 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5931 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5932 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5933 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5934 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5935 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5936 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5937 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5938 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5939 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5940 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5941 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5942 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5943 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5944 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5945 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5946 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5947 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5948 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5949 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5950 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5951 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R616 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M5952 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5953 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5954 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5955 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5956 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5957 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5958 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5959 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R617 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R618 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R619 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M5960 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5961 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5962 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5963 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5964 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5965 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5966 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M5967 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5968 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5969 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5970 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5971 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M5972 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5973 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5974 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5975 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M5976 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5977 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5978 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5979 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5980 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5981 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5982 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5983 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R620 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M5984 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5985 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5986 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M5987 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M5988 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5989 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5990 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M5991 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R621 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R622 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R623 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M5992 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5993 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M5994 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M5995 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M5996 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5997 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M5998 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M5999 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6000 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6001 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6002 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6003 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6004 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6005 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6006 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6007 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R624 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M6008 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6009 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6010 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6011 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6012 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6013 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6014 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6015 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R625 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R626 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R627 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M6016 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6017 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6018 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6019 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6020 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6021 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6022 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6023 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6024 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6025 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6026 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6027 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6028 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6029 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6030 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6031 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6032 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6033 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6034 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6035 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6036 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6037 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6038 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6039 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R628 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M6040 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6041 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6042 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6043 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6044 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6045 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6046 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6047 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R629 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R630 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R631 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M6048 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6049 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6050 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6051 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6052 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6053 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6054 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6055 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6056 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6057 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6058 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6059 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6060 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6061 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6062 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6063 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6064 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6065 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6066 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6067 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6068 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6069 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6070 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6071 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R632 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M6072 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6073 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6074 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6075 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6076 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6077 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6078 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6079 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R633 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R634 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R635 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M6080 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6081 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6082 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6083 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6084 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6085 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6086 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6087 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6088 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6089 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6090 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6091 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6092 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6093 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6094 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6095 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6096 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6097 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6098 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6099 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6100 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6101 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6102 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6103 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R636 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M6104 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6105 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6106 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6107 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6108 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6109 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6110 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6111 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R637 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R638 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R639 9BitDac_0/8BitDac_1/7BitDac_1/R_in7 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M6112 9BitDac_0/8BitDac_1/switchNew_0/a_86_24# D7 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6113 9BitDac_0/8BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6114 9BitDac_0/8BitDac_1/V_out8 9BitDac_0/8BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/V_out7 9BitDac_0/8BitDac_1/7BitDac_0/V_out7 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6115 9BitDac_0/8BitDac_1/7BitDac_0/V_out7 9BitDac_0/8BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/V_out8 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6116 9BitDac_0/8BitDac_1/switchNew_0/a_86_24# D7 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6117 9BitDac_0/8BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6118 9BitDac_0/8BitDac_1/V_out8 9BitDac_0/8BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/V_out7 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6119 9BitDac_0/8BitDac_1/V_out8 9BitDac_0/8BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/V_out7 9BitDac_0/8BitDac_1/V_out8 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6120 9BitDac_0/8BitDac_1/7BitDac_0/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6121 9BitDac_0/8BitDac_1/7BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6122 9BitDac_0/8BitDac_1/7BitDac_0/V_out7 9BitDac_0/8BitDac_1/7BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6123 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 9BitDac_0/8BitDac_1/7BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/V_out7 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6124 9BitDac_0/8BitDac_1/7BitDac_0/switchNew_0/a_86_24# D6 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6125 9BitDac_0/8BitDac_1/7BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6126 9BitDac_0/8BitDac_1/7BitDac_0/V_out7 9BitDac_0/8BitDac_1/7BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6127 9BitDac_0/8BitDac_1/7BitDac_0/V_out7 9BitDac_0/8BitDac_1/7BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 9BitDac_0/8BitDac_1/7BitDac_0/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6128 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6129 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6130 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6131 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6132 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6133 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6134 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6135 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6136 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6137 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6138 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6139 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6140 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6141 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6142 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6143 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6144 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6145 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6146 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6147 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6148 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6149 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6150 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6151 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6152 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6153 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6154 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6155 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6156 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6157 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6158 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_1/R_in7 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6159 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_1/R_in7 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R640 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_1/R_in7 polyResistor w=2 l=62
M6160 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6161 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6162 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6163 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6164 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6165 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6166 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6167 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R641 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R642 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R643 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M6168 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6169 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6170 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6171 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6172 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6173 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6174 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6175 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6176 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6177 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6178 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6179 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6180 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6181 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6182 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6183 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6184 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6185 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6186 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6187 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6188 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6189 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6190 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6191 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R644 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M6192 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6193 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6194 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6195 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6196 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6197 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6198 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6199 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R645 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R646 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R647 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M6200 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6201 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6202 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6203 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6204 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6205 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6206 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6207 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6208 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6209 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6210 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6211 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6212 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6213 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6214 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6215 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6216 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6217 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6218 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6219 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6220 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6221 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6222 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6223 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R648 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M6224 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6225 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6226 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6227 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6228 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6229 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6230 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6231 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R649 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R650 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R651 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M6232 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6233 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6234 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6235 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6236 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6237 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6238 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6239 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6240 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6241 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6242 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6243 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6244 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6245 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6246 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6247 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6248 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6249 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6250 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6251 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6252 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6253 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6254 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6255 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R652 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M6256 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6257 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6258 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6259 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6260 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6261 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6262 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6263 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R653 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R654 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R655 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M6264 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6265 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6266 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6267 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6268 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6269 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6270 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6271 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6272 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6273 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6274 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6275 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6276 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6277 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6278 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6279 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R656 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M6280 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6281 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6282 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6283 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6284 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6285 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6286 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6287 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R657 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R658 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R659 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M6288 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6289 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6290 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6291 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6292 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6293 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6294 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6295 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6296 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6297 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6298 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6299 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6300 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6301 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6302 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6303 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6304 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6305 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6306 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6307 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6308 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6309 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6310 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6311 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R660 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M6312 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6313 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6314 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6315 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6316 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6317 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6318 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6319 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R661 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R662 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R663 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M6320 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6321 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6322 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6323 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6324 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6325 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6326 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6327 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6328 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6329 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6330 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6331 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6332 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6333 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6334 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6335 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6336 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6337 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6338 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6339 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6340 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6341 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6342 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6343 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R664 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M6344 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6345 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6346 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6347 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6348 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6349 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6350 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6351 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R665 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R666 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R667 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M6352 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6353 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6354 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6355 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6356 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6357 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6358 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6359 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6360 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6361 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6362 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6363 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6364 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6365 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6366 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6367 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6368 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6369 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6370 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6371 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6372 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6373 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6374 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6375 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R668 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M6376 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6377 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6378 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6379 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6380 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6381 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6382 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6383 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R669 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R670 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R671 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M6384 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6385 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6386 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6387 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6388 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6389 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6390 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6391 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6392 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6393 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6394 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6395 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6396 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6397 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6398 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6399 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6400 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6401 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6402 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6403 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6404 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6405 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6406 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6407 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R672 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M6408 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6409 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6410 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6411 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6412 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6413 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6414 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6415 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R673 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R674 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R675 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M6416 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6417 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6418 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6419 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6420 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6421 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6422 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6423 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6424 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6425 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6426 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6427 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6428 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6429 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6430 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6431 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6432 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6433 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6434 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6435 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6436 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6437 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6438 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6439 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R676 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M6440 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6441 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6442 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6443 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6444 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6445 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6446 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6447 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R677 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R678 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R679 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M6448 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6449 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6450 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6451 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6452 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6453 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6454 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6455 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6456 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6457 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6458 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6459 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6460 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6461 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6462 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6463 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6464 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6465 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6466 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6467 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6468 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6469 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6470 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6471 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R680 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M6472 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6473 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6474 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6475 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6476 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6477 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6478 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6479 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R681 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R682 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R683 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M6480 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6481 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6482 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6483 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6484 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6485 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6486 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6487 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6488 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6489 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6490 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6491 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6492 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6493 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6494 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6495 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6496 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6497 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6498 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6499 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6500 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6501 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6502 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6503 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R684 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M6504 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6505 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6506 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6507 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6508 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6509 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6510 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6511 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R685 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R686 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R687 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M6512 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6513 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6514 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6515 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6516 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6517 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6518 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6519 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6520 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6521 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6522 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6523 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6524 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6525 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6526 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6527 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R688 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M6528 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6529 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6530 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6531 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6532 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6533 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6534 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6535 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R689 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R690 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R691 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M6536 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6537 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6538 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6539 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6540 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6541 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6542 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6543 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6544 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6545 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6546 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6547 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6548 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6549 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6550 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6551 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6552 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6553 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6554 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6555 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6556 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6557 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6558 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6559 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R692 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M6560 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6561 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6562 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6563 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6564 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6565 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6566 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6567 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R693 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R694 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R695 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M6568 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6569 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6570 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6571 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6572 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6573 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6574 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6575 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6576 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6577 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6578 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6579 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6580 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6581 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6582 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6583 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6584 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6585 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6586 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6587 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6588 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6589 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6590 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6591 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R696 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M6592 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6593 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6594 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6595 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6596 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6597 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6598 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6599 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R697 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R698 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R699 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M6600 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6601 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6602 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6603 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6604 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6605 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6606 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6607 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6608 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6609 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6610 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6611 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6612 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6613 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6614 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6615 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6616 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6617 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6618 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6619 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6620 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6621 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6622 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6623 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R700 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M6624 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6625 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6626 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6627 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6628 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6629 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6630 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6631 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R701 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R702 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R703 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/R_in6 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M6632 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6633 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6634 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6635 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6636 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6637 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6638 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6639 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6640 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6641 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6642 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6643 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6644 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6645 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6646 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6647 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6648 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6649 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6650 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6651 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6652 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6653 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6654 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6655 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6656 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6657 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6658 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6659 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6660 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6661 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6662 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/R_in6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6663 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/R_in6 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R704 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/R_in6 polyResistor w=2 l=62
M6664 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6665 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6666 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6667 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6668 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6669 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6670 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6671 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R705 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R706 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R707 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M6672 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6673 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6674 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6675 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6676 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6677 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6678 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6679 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6680 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6681 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6682 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6683 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6684 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6685 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6686 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6687 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6688 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6689 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6690 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6691 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6692 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6693 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6694 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6695 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R708 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M6696 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6697 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6698 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6699 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6700 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6701 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6702 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6703 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R709 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R710 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R711 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M6704 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6705 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6706 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6707 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6708 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6709 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6710 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6711 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6712 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6713 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6714 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6715 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6716 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6717 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6718 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6719 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6720 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6721 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6722 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6723 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6724 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6725 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6726 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6727 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R712 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M6728 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6729 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6730 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6731 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6732 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6733 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6734 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6735 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R713 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R714 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R715 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M6736 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6737 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6738 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6739 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6740 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6741 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6742 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6743 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6744 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6745 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6746 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6747 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6748 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6749 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6750 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6751 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6752 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6753 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6754 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6755 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6756 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6757 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6758 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6759 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R716 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M6760 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6761 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6762 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6763 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6764 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6765 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6766 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6767 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R717 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R718 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R719 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M6768 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6769 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6770 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6771 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6772 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6773 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6774 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6775 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6776 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6777 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6778 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6779 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6780 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6781 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6782 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6783 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R720 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M6784 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6785 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6786 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6787 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6788 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6789 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6790 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6791 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R721 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R722 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R723 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M6792 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6793 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6794 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6795 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6796 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6797 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6798 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6799 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6800 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6801 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6802 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6803 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6804 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6805 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6806 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6807 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6808 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6809 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6810 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6811 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6812 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6813 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6814 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6815 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R724 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M6816 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6817 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6818 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6819 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6820 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6821 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6822 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6823 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R725 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R726 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R727 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M6824 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6825 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6826 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6827 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6828 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6829 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6830 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6831 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6832 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6833 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6834 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6835 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6836 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6837 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6838 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6839 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6840 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6841 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6842 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6843 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6844 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6845 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6846 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6847 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R728 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M6848 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6849 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6850 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6851 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6852 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6853 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6854 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6855 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R729 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R730 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R731 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M6856 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6857 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6858 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6859 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6860 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6861 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6862 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6863 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6864 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6865 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6866 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6867 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6868 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6869 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6870 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6871 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6872 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6873 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6874 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6875 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6876 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6877 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6878 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6879 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R732 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M6880 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6881 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6882 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6883 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6884 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6885 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6886 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6887 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R733 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R734 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R735 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M6888 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6889 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6890 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6891 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6892 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6893 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6894 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6895 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6896 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6897 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6898 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6899 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6900 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6901 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6902 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6903 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6904 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6905 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6906 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6907 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6908 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6909 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6910 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6911 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R736 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M6912 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6913 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6914 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6915 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6916 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6917 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6918 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6919 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R737 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R738 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R739 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M6920 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6921 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6922 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6923 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6924 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6925 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6926 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6927 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6928 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6929 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6930 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6931 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6932 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6933 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6934 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6935 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6936 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6937 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6938 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6939 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6940 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6941 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6942 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6943 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R740 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M6944 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6945 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6946 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6947 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6948 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6949 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6950 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6951 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R741 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R742 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R743 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M6952 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6953 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6954 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6955 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6956 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6957 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6958 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6959 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6960 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6961 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6962 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M6963 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M6964 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6965 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6966 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6967 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6968 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6969 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6970 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6971 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6972 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6973 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6974 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6975 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R744 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M6976 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6977 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6978 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M6979 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M6980 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6981 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6982 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M6983 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R745 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R746 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R747 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M6984 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6985 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6986 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6987 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6988 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6989 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6990 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M6991 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6992 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6993 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M6994 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M6995 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M6996 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6997 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M6998 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M6999 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7000 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7001 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7002 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7003 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7004 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7005 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7006 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7007 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R748 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M7008 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7009 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7010 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7011 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7012 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7013 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7014 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7015 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R749 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R750 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R751 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M7016 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7017 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7018 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7019 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7020 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7021 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7022 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7023 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7024 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7025 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7026 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7027 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7028 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7029 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7030 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7031 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R752 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M7032 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7033 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7034 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7035 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7036 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7037 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7038 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7039 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R753 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R754 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R755 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M7040 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7041 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7042 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7043 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7044 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7045 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7046 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7047 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7048 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7049 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7050 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7051 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7052 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7053 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7054 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7055 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7056 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7057 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7058 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7059 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7060 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7061 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7062 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7063 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R756 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M7064 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7065 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7066 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7067 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7068 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7069 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7070 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7071 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R757 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R758 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R759 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M7072 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7073 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7074 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7075 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7076 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7077 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7078 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7079 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7080 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7081 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7082 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7083 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7084 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7085 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7086 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7087 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7088 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7089 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7090 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7091 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7092 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7093 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7094 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7095 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R760 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M7096 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7097 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7098 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7099 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7100 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7101 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7102 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7103 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R761 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R762 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R763 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M7104 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7105 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7106 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7107 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7108 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7109 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7110 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7111 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7112 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7113 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7114 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7115 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7116 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7117 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7118 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7119 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7120 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7121 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7122 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7123 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7124 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7125 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7126 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7127 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R764 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M7128 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7129 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7130 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7131 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7132 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7133 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7134 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7135 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R765 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R766 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R767 9BitDac_0/8BitDac_1/R_in8 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M7136 9BitDac_0/switchNew_0/a_86_24# D8 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7137 9BitDac_0/switchNew_0/a_105_21# 9BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7138 9BitDac_0/V_out9 9BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/V_out8 9BitDac_0/8BitDac_0/V_out8 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7139 9BitDac_0/8BitDac_0/V_out8 9BitDac_0/switchNew_0/a_105_21# 9BitDac_0/V_out9 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7140 9BitDac_0/switchNew_0/a_86_24# D8 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7141 9BitDac_0/switchNew_0/a_105_21# 9BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7142 9BitDac_0/V_out9 9BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_1/V_out8 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7143 9BitDac_0/V_out9 9BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_1/V_out8 9BitDac_0/V_out9 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7144 9BitDac_0/8BitDac_0/7BitDac_1/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7145 9BitDac_0/8BitDac_0/7BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7146 9BitDac_0/8BitDac_0/7BitDac_1/V_out7 9BitDac_0/8BitDac_0/7BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7147 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 9BitDac_0/8BitDac_0/7BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/V_out7 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7148 9BitDac_0/8BitDac_0/7BitDac_1/switchNew_0/a_86_24# D6 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7149 9BitDac_0/8BitDac_0/7BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7150 9BitDac_0/8BitDac_0/7BitDac_1/V_out7 9BitDac_0/8BitDac_0/7BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7151 9BitDac_0/8BitDac_0/7BitDac_1/V_out7 9BitDac_0/8BitDac_0/7BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 9BitDac_0/8BitDac_0/7BitDac_1/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7152 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7153 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7154 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7155 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7156 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7157 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7158 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7159 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7160 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7161 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7162 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7163 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7164 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7165 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7166 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7167 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7168 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7169 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7170 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7171 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7172 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7173 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7174 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7175 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7176 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7177 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7178 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7179 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7180 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7181 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7182 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_1/R_in8 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7183 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_1/R_in8 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R768 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_1/R_in8 polyResistor w=2 l=62
M7184 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7185 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7186 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7187 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7188 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7189 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7190 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7191 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R769 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R770 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R771 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M7192 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7193 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7194 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7195 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7196 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7197 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7198 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7199 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7200 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7201 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7202 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7203 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7204 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7205 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7206 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7207 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7208 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7209 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7210 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7211 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7212 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7213 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7214 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7215 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R772 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M7216 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7217 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7218 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7219 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7220 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7221 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7222 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7223 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R773 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R774 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R775 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M7224 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7225 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7226 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7227 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7228 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7229 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7230 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7231 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7232 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7233 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7234 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7235 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7236 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7237 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7238 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7239 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7240 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7241 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7242 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7243 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7244 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7245 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7246 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7247 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R776 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M7248 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7249 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7250 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7251 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7252 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7253 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7254 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7255 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R777 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R778 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R779 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M7256 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7257 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7258 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7259 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7260 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7261 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7262 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7263 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7264 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7265 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7266 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7267 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7268 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7269 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7270 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7271 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7272 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7273 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7274 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7275 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7276 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7277 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7278 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7279 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R780 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M7280 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7281 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7282 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7283 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7284 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7285 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7286 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7287 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R781 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R782 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R783 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M7288 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7289 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7290 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7291 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7292 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7293 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7294 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7295 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7296 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7297 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7298 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7299 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7300 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7301 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7302 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7303 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R784 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M7304 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7305 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7306 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7307 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7308 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7309 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7310 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7311 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R785 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R786 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R787 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M7312 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7313 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7314 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7315 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7316 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7317 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7318 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7319 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7320 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7321 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7322 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7323 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7324 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7325 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7326 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7327 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7328 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7329 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7330 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7331 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7332 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7333 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7334 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7335 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R788 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M7336 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7337 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7338 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7339 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7340 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7341 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7342 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7343 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R789 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R790 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R791 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M7344 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7345 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7346 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7347 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7348 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7349 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7350 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7351 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7352 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7353 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7354 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7355 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7356 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7357 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7358 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7359 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7360 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7361 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7362 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7363 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7364 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7365 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7366 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7367 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R792 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M7368 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7369 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7370 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7371 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7372 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7373 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7374 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7375 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R793 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R794 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R795 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M7376 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7377 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7378 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7379 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7380 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7381 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7382 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7383 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7384 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7385 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7386 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7387 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7388 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7389 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7390 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7391 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7392 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7393 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7394 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7395 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7396 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7397 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7398 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7399 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R796 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M7400 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7401 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7402 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7403 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7404 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7405 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7406 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7407 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R797 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R798 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R799 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M7408 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7409 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7410 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7411 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7412 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7413 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7414 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7415 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7416 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7417 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7418 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7419 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7420 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7421 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7422 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7423 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7424 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7425 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7426 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7427 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7428 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7429 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7430 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7431 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R800 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M7432 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7433 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7434 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7435 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7436 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7437 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7438 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7439 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R801 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R802 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R803 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M7440 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7441 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7442 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7443 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7444 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7445 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7446 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7447 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7448 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7449 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7450 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7451 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7452 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7453 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7454 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7455 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7456 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7457 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7458 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7459 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7460 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7461 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7462 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7463 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R804 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M7464 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7465 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7466 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7467 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7468 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7469 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7470 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7471 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R805 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R806 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R807 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M7472 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7473 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7474 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7475 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7476 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7477 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7478 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7479 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7480 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7481 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7482 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7483 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7484 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7485 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7486 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7487 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7488 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7489 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7490 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7491 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7492 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7493 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7494 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7495 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R808 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M7496 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7497 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7498 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7499 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7500 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7501 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7502 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7503 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R809 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R810 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R811 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M7504 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7505 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7506 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7507 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7508 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7509 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7510 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7511 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7512 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7513 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7514 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7515 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7516 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7517 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7518 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7519 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7520 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7521 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7522 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7523 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7524 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7525 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7526 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7527 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R812 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M7528 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7529 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7530 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7531 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7532 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7533 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7534 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7535 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R813 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R814 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R815 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M7536 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7537 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7538 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7539 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7540 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7541 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7542 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7543 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7544 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7545 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7546 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7547 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7548 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7549 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7550 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7551 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R816 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M7552 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7553 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7554 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7555 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7556 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7557 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7558 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7559 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R817 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R818 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R819 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M7560 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7561 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7562 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7563 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7564 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7565 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7566 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7567 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7568 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7569 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7570 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7571 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7572 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7573 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7574 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7575 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7576 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7577 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7578 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7579 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7580 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7581 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7582 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7583 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R820 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M7584 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7585 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7586 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7587 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7588 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7589 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7590 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7591 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R821 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R822 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R823 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M7592 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7593 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7594 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7595 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7596 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7597 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7598 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7599 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7600 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7601 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7602 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7603 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7604 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7605 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7606 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7607 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7608 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7609 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7610 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7611 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7612 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7613 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7614 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7615 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R824 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M7616 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7617 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7618 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7619 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7620 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7621 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7622 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7623 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R825 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R826 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R827 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M7624 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7625 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7626 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7627 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7628 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7629 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7630 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7631 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7632 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7633 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7634 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7635 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7636 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7637 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7638 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7639 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7640 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7641 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7642 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7643 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7644 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7645 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7646 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7647 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R828 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M7648 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7649 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7650 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7651 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7652 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7653 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7654 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7655 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R829 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R830 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R831 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/R_in6 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M7656 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7657 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7658 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7659 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7660 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7661 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7662 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7663 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7664 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7665 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7666 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7667 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7668 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7669 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7670 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7671 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7672 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7673 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7674 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7675 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7676 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7677 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7678 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7679 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7680 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7681 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7682 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7683 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7684 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7685 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7686 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/R_in6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7687 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/R_in6 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R832 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/R_in6 polyResistor w=2 l=62
M7688 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7689 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7690 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7691 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7692 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7693 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7694 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7695 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R833 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R834 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R835 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M7696 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7697 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7698 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7699 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7700 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7701 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7702 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7703 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7704 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7705 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7706 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7707 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7708 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7709 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7710 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7711 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7712 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7713 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7714 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7715 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7716 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7717 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7718 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7719 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R836 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M7720 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7721 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7722 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7723 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7724 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7725 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7726 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7727 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R837 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R838 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R839 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M7728 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7729 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7730 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7731 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7732 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7733 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7734 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7735 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7736 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7737 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7738 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7739 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7740 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7741 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7742 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7743 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7744 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7745 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7746 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7747 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7748 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7749 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7750 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7751 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R840 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M7752 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7753 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7754 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7755 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7756 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7757 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7758 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7759 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R841 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R842 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R843 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M7760 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7761 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7762 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7763 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7764 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7765 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7766 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7767 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7768 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7769 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7770 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7771 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7772 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7773 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7774 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7775 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7776 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7777 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7778 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7779 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7780 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7781 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7782 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7783 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R844 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M7784 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7785 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7786 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7787 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7788 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7789 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7790 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7791 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R845 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R846 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R847 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M7792 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7793 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7794 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7795 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7796 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7797 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7798 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7799 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7800 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7801 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7802 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7803 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7804 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7805 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7806 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7807 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R848 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M7808 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7809 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7810 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7811 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7812 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7813 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7814 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7815 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R849 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R850 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R851 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M7816 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7817 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7818 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7819 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7820 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7821 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7822 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7823 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7824 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7825 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7826 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7827 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7828 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7829 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7830 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7831 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7832 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7833 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7834 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7835 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7836 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7837 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7838 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7839 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R852 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M7840 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7841 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7842 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7843 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7844 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7845 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7846 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7847 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R853 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R854 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R855 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M7848 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7849 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7850 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7851 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7852 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7853 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7854 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7855 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7856 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7857 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7858 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7859 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7860 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7861 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7862 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7863 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7864 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7865 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7866 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7867 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7868 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7869 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7870 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7871 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R856 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M7872 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7873 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7874 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7875 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7876 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7877 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7878 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7879 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R857 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R858 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R859 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M7880 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7881 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7882 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7883 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7884 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7885 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7886 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7887 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7888 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7889 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7890 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7891 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7892 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7893 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7894 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7895 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7896 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7897 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7898 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7899 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7900 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7901 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7902 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7903 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R860 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M7904 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7905 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7906 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7907 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7908 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7909 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7910 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7911 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R861 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R862 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R863 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M7912 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7913 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7914 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7915 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7916 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7917 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7918 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7919 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7920 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7921 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7922 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7923 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7924 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7925 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7926 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7927 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7928 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7929 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7930 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7931 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7932 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7933 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7934 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7935 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R864 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M7936 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7937 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7938 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7939 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7940 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7941 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7942 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7943 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R865 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R866 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R867 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M7944 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7945 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7946 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7947 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7948 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7949 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7950 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7951 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7952 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7953 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7954 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7955 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7956 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7957 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7958 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7959 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7960 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7961 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7962 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7963 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7964 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7965 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7966 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7967 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R868 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M7968 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7969 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7970 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7971 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7972 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7973 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7974 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7975 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R869 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R870 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R871 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M7976 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7977 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7978 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7979 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M7980 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7981 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7982 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M7983 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7984 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7985 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7986 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M7987 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M7988 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7989 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7990 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M7991 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M7992 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7993 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M7994 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M7995 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M7996 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7997 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M7998 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M7999 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R872 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M8000 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8001 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8002 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8003 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8004 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8005 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8006 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8007 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R873 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R874 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R875 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M8008 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8009 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8010 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8011 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8012 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8013 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8014 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8015 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8016 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8017 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8018 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8019 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8020 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8021 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8022 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8023 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8024 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8025 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8026 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8027 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8028 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8029 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8030 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8031 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R876 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M8032 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8033 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8034 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8035 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8036 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8037 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8038 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8039 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R877 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R878 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R879 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M8040 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8041 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8042 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8043 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8044 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8045 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8046 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8047 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8048 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8049 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8050 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8051 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8052 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8053 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8054 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8055 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R880 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M8056 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8057 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8058 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8059 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8060 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8061 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8062 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8063 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R881 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R882 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R883 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M8064 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8065 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8066 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8067 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8068 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8069 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8070 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8071 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8072 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8073 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8074 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8075 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8076 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8077 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8078 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8079 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8080 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8081 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8082 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8083 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8084 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8085 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8086 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8087 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R884 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M8088 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8089 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8090 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8091 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8092 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8093 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8094 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8095 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R885 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R886 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R887 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M8096 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8097 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8098 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8099 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8100 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8101 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8102 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8103 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8104 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8105 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8106 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8107 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8108 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8109 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8110 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8111 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8112 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8113 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8114 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8115 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8116 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8117 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8118 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8119 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R888 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M8120 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8121 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8122 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8123 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8124 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8125 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8126 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8127 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R889 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R890 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R891 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M8128 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8129 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8130 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8131 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8132 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8133 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8134 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8135 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8136 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8137 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8138 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8139 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8140 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8141 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8142 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8143 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8144 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8145 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8146 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8147 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8148 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8149 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8150 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8151 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R892 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M8152 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8153 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8154 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8155 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8156 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8157 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8158 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8159 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R893 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R894 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R895 9BitDac_0/8BitDac_0/7BitDac_1/R_in7 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M8160 9BitDac_0/8BitDac_0/switchNew_0/a_86_24# D7 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8161 9BitDac_0/8BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8162 9BitDac_0/8BitDac_0/V_out8 9BitDac_0/8BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/V_out7 9BitDac_0/8BitDac_0/7BitDac_0/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8163 9BitDac_0/8BitDac_0/7BitDac_0/V_out7 9BitDac_0/8BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/V_out8 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8164 9BitDac_0/8BitDac_0/switchNew_0/a_86_24# D7 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8165 9BitDac_0/8BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8166 9BitDac_0/8BitDac_0/V_out8 9BitDac_0/8BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/V_out7 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8167 9BitDac_0/8BitDac_0/V_out8 9BitDac_0/8BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/V_out7 9BitDac_0/8BitDac_0/V_out8 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8168 9BitDac_0/8BitDac_0/7BitDac_0/switchNew_0/a_86_24# D6 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8169 9BitDac_0/8BitDac_0/7BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8170 9BitDac_0/8BitDac_0/7BitDac_0/V_out7 9BitDac_0/8BitDac_0/7BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8171 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 9BitDac_0/8BitDac_0/7BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/V_out7 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8172 9BitDac_0/8BitDac_0/7BitDac_0/switchNew_0/a_86_24# D6 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8173 9BitDac_0/8BitDac_0/7BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8174 9BitDac_0/8BitDac_0/7BitDac_0/V_out7 9BitDac_0/8BitDac_0/7BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8175 9BitDac_0/8BitDac_0/7BitDac_0/V_out7 9BitDac_0/8BitDac_0/7BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 9BitDac_0/8BitDac_0/7BitDac_0/V_out7 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8176 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8177 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8178 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8179 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8180 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8181 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8182 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8183 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8184 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8185 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8186 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8187 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8188 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8189 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8190 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8191 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8192 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8193 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8194 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8195 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8196 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8197 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8198 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8199 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8200 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8201 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8202 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8203 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8204 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8205 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8206 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_1/R_in7 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8207 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_1/R_in7 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R896 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_1/R_in7 polyResistor w=2 l=62
M8208 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8209 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8210 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8211 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8212 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8213 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8214 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8215 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R897 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R898 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R899 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M8216 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8217 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8218 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8219 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8220 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8221 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8222 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8223 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8224 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8225 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8226 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8227 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8228 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8229 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8230 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8231 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8232 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8233 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8234 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8235 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8236 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8237 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8238 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8239 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R900 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M8240 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8241 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8242 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8243 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8244 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8245 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8246 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8247 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R901 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R902 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R903 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M8248 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8249 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8250 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8251 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8252 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8253 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8254 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8255 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8256 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8257 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8258 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8259 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8260 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8261 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8262 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8263 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8264 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8265 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8266 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8267 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8268 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8269 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8270 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8271 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R904 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M8272 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8273 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8274 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8275 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8276 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8277 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8278 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8279 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R905 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R906 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R907 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M8280 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8281 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8282 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8283 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8284 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8285 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8286 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8287 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8288 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8289 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8290 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8291 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8292 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8293 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8294 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8295 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8296 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8297 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8298 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8299 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8300 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8301 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8302 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8303 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R908 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M8304 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8305 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8306 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8307 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8308 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8309 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8310 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8311 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R909 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R910 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R911 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M8312 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8313 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8314 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8315 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8316 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8317 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8318 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8319 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8320 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8321 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8322 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8323 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8324 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8325 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8326 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8327 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R912 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M8328 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8329 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8330 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8331 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8332 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8333 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8334 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8335 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R913 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R914 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R915 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M8336 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8337 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8338 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8339 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8340 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8341 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8342 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8343 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8344 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8345 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8346 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8347 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8348 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8349 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8350 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8351 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8352 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8353 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8354 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8355 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8356 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8357 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8358 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8359 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R916 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M8360 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8361 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8362 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8363 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8364 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8365 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8366 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8367 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R917 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R918 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R919 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M8368 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8369 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8370 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8371 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8372 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8373 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8374 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8375 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8376 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8377 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8378 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8379 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8380 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8381 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8382 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8383 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8384 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8385 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8386 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8387 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8388 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8389 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8390 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8391 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R920 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M8392 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8393 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8394 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8395 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8396 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8397 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8398 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8399 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R921 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R922 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R923 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M8400 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8401 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8402 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8403 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8404 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8405 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8406 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8407 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8408 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8409 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8410 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8411 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8412 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8413 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8414 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8415 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8416 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8417 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8418 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8419 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8420 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8421 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8422 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8423 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R924 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M8424 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8425 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8426 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8427 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8428 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8429 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8430 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8431 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R925 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R926 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R927 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M8432 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8433 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8434 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8435 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8436 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8437 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8438 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8439 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8440 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8441 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8442 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8443 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8444 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8445 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8446 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8447 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8448 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8449 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8450 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8451 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8452 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8453 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8454 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8455 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R928 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/R_in5 polyResistor w=2 l=62
M8456 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8457 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8458 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8459 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8460 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8461 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8462 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8463 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R929 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R930 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R931 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M8464 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8465 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8466 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8467 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8468 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8469 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8470 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8471 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8472 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8473 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8474 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8475 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8476 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8477 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8478 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8479 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8480 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8481 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8482 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8483 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8484 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8485 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8486 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8487 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R932 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M8488 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8489 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8490 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8491 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8492 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8493 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8494 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8495 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R933 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R934 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R935 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M8496 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8497 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8498 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8499 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8500 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8501 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8502 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8503 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8504 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8505 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8506 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8507 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8508 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8509 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8510 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8511 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8512 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8513 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8514 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8515 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8516 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8517 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8518 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8519 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R936 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M8520 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8521 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8522 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8523 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8524 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8525 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8526 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8527 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R937 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R938 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R939 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M8528 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8529 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8530 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8531 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8532 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8533 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8534 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8535 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8536 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8537 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8538 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8539 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8540 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8541 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8542 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8543 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8544 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8545 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8546 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8547 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8548 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8549 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8550 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8551 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R940 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M8552 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8553 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8554 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8555 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8556 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8557 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8558 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8559 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R941 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R942 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R943 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M8560 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8561 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8562 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8563 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8564 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8565 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8566 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8567 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8568 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8569 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8570 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8571 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8572 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8573 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8574 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8575 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R944 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M8576 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8577 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8578 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8579 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8580 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8581 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8582 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8583 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R945 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R946 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R947 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M8584 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8585 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8586 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8587 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8588 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8589 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8590 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8591 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8592 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8593 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8594 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8595 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8596 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8597 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8598 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8599 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8600 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8601 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8602 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8603 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8604 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8605 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8606 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8607 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R948 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M8608 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8609 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8610 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8611 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8612 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8613 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8614 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8615 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R949 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R950 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R951 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M8616 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8617 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8618 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8619 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8620 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8621 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8622 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8623 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8624 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8625 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8626 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8627 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8628 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8629 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8630 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8631 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8632 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8633 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8634 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8635 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8636 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8637 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8638 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8639 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R952 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M8640 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8641 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8642 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8643 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8644 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8645 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8646 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8647 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R953 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R954 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R955 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M8648 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8649 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8650 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8651 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8652 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8653 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8654 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8655 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8656 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8657 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8658 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8659 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8660 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8661 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8662 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8663 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8664 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8665 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8666 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8667 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8668 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8669 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8670 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8671 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R956 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M8672 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8673 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8674 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8675 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8676 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8677 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8678 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8679 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R957 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R958 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R959 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/R_in6 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M8680 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8681 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8682 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8683 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8684 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# D5 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8685 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8686 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8687 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8688 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8689 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8690 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8691 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8692 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8693 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8694 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8695 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8696 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8697 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8698 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8699 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8700 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8701 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8702 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8703 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8704 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8705 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8706 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8707 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8708 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8709 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8710 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/R_in6 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8711 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/R_in6 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R960 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/R_in6 polyResistor w=2 l=62
M8712 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8713 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8714 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8715 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8716 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8717 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8718 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8719 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R961 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R962 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R963 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M8720 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8721 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8722 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8723 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8724 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8725 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8726 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8727 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8728 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8729 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8730 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8731 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8732 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8733 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8734 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8735 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8736 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8737 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8738 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8739 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8740 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8741 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8742 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8743 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R964 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M8744 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8745 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8746 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8747 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8748 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8749 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8750 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8751 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R965 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R966 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R967 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M8752 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8753 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8754 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8755 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8756 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8757 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8758 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8759 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8760 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8761 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8762 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8763 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8764 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8765 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8766 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8767 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8768 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8769 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8770 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8771 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8772 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8773 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8774 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8775 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R968 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M8776 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8777 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8778 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8779 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8780 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8781 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8782 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8783 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R969 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R970 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R971 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M8784 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8785 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8786 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8787 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8788 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8789 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8790 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8791 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8792 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8793 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8794 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8795 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8796 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8797 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8798 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8799 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8800 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8801 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8802 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8803 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8804 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8805 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8806 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8807 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R972 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M8808 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8809 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8810 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8811 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8812 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8813 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8814 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8815 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R973 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R974 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R975 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M8816 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8817 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8818 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8819 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8820 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8821 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8822 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8823 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8824 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8825 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8826 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8827 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8828 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8829 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8830 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8831 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R976 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/R_in4 polyResistor w=2 l=62
M8832 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8833 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8834 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8835 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8836 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8837 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8838 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8839 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R977 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R978 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R979 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M8840 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8841 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8842 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8843 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8844 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8845 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8846 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8847 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8848 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8849 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8850 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8851 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8852 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8853 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8854 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8855 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8856 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8857 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8858 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8859 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8860 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8861 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8862 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8863 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R980 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M8864 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8865 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8866 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8867 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8868 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8869 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8870 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8871 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R981 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R982 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R983 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M8872 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8873 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8874 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8875 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8876 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8877 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8878 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8879 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8880 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8881 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8882 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8883 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8884 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8885 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8886 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8887 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8888 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8889 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8890 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8891 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8892 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8893 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8894 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8895 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R984 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M8896 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8897 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8898 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8899 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8900 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8901 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8902 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8903 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R985 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R986 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R987 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M8904 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8905 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8906 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8907 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8908 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8909 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8910 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8911 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8912 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8913 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8914 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8915 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8916 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8917 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8918 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8919 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8920 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8921 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8922 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8923 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8924 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8925 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8926 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8927 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R988 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M8928 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8929 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8930 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8931 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8932 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8933 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8934 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8935 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R989 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R990 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R991 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M8936 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8937 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8938 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8939 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8940 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# D4 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8941 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8942 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8943 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/V_out5 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8944 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8945 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8946 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8947 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8948 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8949 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8950 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8951 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8952 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8953 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8954 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8955 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8956 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8957 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8958 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8959 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R992 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/R_in5 polyResistor w=2 l=62
M8960 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8961 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8962 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8963 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8964 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8965 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8966 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8967 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R993 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R994 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R995 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M8968 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8969 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8970 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M8971 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M8972 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8973 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8974 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M8975 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8976 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8977 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8978 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8979 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M8980 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8981 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8982 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M8983 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M8984 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8985 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8986 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8987 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8988 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8989 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8990 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8991 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R996 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M8992 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8993 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M8994 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M8995 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M8996 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8997 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M8998 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M8999 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R997 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R998 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R999 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M9000 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9001 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9002 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M9003 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M9004 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9005 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9006 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M9007 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9008 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9009 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9010 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M9011 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M9012 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9013 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9014 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M9015 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M9016 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9017 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9018 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M9019 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M9020 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9021 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9022 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M9023 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1000 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/R_in3 polyResistor w=2 l=62
M9024 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9025 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9026 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M9027 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M9028 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9029 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9030 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M9031 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1001 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R1002 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R1003 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M9032 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9033 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9034 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M9035 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M9036 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9037 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9038 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M9039 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9040 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9041 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9042 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M9043 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M9044 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9045 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9046 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M9047 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M9048 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9049 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9050 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M9051 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M9052 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9053 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9054 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M9055 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1004 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M9056 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9057 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9058 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M9059 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M9060 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9061 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9062 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M9063 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1005 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R1006 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R1007 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
M9064 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9065 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9066 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M9067 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M9068 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9069 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9070 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M9071 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M9072 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9073 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9074 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M9075 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M9076 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9077 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9078 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M9079 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1008 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/R_in4 polyResistor w=2 l=62
M9080 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9081 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9082 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M9083 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M9084 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9085 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9086 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M9087 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1009 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/gamma polyResistor w=2 l=62
R1010 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/beta polyResistor w=2 l=62
R1011 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/alpha polyResistor w=2 l=62
M9088 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9089 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9090 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M9091 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M9092 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9093 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9094 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M9095 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9096 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9097 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9098 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M9099 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M9100 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9101 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9102 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M9103 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M9104 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9105 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9106 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M9107 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M9108 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9109 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9110 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M9111 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1012 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/delta polyResistor w=2 l=62
M9112 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9113 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9114 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M9115 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M9116 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9117 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9118 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M9119 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1013 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/gamma polyResistor w=2 l=62
R1014 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/beta polyResistor w=2 l=62
R1015 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/alpha polyResistor w=2 l=62
M9120 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9121 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9122 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M9123 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M9124 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# D3 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9125 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9126 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M9127 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9128 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9129 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9130 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=210 pd=102 as=210 ps=102
M9131 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=121 ps=88
M9132 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9133 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9134 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M9135 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M9136 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9137 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9138 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M9139 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M9140 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9141 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9142 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M9143 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1016 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/R_in3 polyResistor w=2 l=62
M9144 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9145 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9146 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M9147 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M9148 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9149 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9150 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M9151 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1017 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/gamma polyResistor w=2 l=62
R1018 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/beta polyResistor w=2 l=62
R1019 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/alpha polyResistor w=2 l=62
M9152 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9153 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9154 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M9155 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M9156 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# D2 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9157 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9158 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
M9159 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9160 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9161 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9162 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M9163 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd nfet w=5 l=2
+  ad=137 pd=104 as=0 ps=0
M9164 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# D1 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9165 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9166 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=0 pd=0 as=121 ps=88
M9167 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_2/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 pfet w=10 l=2
+  ad=0 pd=0 as=210 ps=102
M9168 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9169 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9170 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M9171 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M9172 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9173 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9174 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M9175 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_1/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_198_n130# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1020 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/delta polyResistor w=2 l=62
M9176 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9177 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# VA VA pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M9178 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
M9179 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# gnd nfet w=5 l=2
+  ad=51 pd=40 as=0 ps=0
M9180 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# D0 gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9181 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# gnd gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M9182 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_86_24# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta gnd nfet w=5 l=2
+  ad=0 pd=0 as=35 ps=24
M9183 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/switchNew_0/a_105_21# 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/m1_201_n40# pfet w=10 l=2
+  ad=0 pd=0 as=70 ps=34
R1021 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/gamma polyResistor w=2 l=62
R1022 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/beta polyResistor w=2 l=62
R1023 R_in10 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/alpha polyResistor w=2 l=62
C1 D6 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 5.36fF
C2 VA D5 2.83fF
C3 D4 VA 7.03fF
C4 D6 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 5.31fF
C5 D6 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/V_out6 5.31fF
C6 D0 VA 41.71fF
C7 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/V_out6 D6 5.31fF
C8 D6 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 5.31fF
C9 D2 D3 3.38fF
C10 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/V_out6 D6 5.31fF
C11 D2 VA 45.52fF
C12 D2 D1 233.09fF
C13 D3 VA 63.18fF
C14 D3 D1 44.63fF
C15 D1 VA 122.26fF
C16 D2 9BitDac_0/8BitDac_0/7BitDac_0/V_out7 3.39fF
C17 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 D6 5.31fF
C18 D6 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/V_out6 5.31fF
C19 9BitDac_1/8BitDac_0/7BitDac_0/V_out7 D2 3.39fF
C20 D5 gnd 5.22fF
C21 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C22 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C23 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C24 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C25 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C26 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C27 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C28 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C29 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C30 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C31 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C32 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C33 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C34 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C35 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C36 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C37 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C38 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C39 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C40 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C41 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C42 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C43 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C44 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C45 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C46 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C47 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C48 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C49 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C50 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C51 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C52 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C53 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C54 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C55 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C56 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C57 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C58 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C59 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C60 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C61 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C62 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C63 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C64 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C65 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C66 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C67 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C68 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C69 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C70 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C71 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C72 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C73 9BitDac_0/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 gnd 2.06fF
C74 9BitDac_0/8BitDac_0/7BitDac_1/V_out7 gnd 2.40fF
C75 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C76 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C77 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C78 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C79 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C80 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C81 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C82 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C83 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C84 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C85 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C86 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C87 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C88 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C89 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C90 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C91 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C92 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C93 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C94 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C95 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C96 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C97 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C98 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C99 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C100 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C101 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C102 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C103 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C104 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C105 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C106 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C107 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C108 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C109 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C110 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C111 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C112 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C113 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C114 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C115 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C116 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C117 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C118 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C119 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C120 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C121 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C122 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C123 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C124 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C125 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C126 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C127 9BitDac_0/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 gnd 2.06fF
C128 9BitDac_0/8BitDac_1/V_out8 gnd 2.32fF
C129 9BitDac_0/8BitDac_0/V_out8 gnd 2.04fF
C130 VA gnd 1849.19fF
C131 9BitDac_0/8BitDac_1/R_in8 gnd 2.05fF
C132 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C133 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C134 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C135 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C136 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C137 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C138 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C139 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C140 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C141 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C142 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C143 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C144 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C145 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C146 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C147 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C148 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C149 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C150 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C151 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C152 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C153 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C154 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C155 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C156 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C157 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C158 D1 gnd 154.87fF
C159 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C160 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C161 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C162 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C163 D3 gnd 3.53fF
C164 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C165 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C166 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C167 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C168 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C169 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C170 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C171 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C172 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C173 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C174 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C175 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C176 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C177 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C178 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C179 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C180 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C181 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C182 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C183 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C184 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C185 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C186 9BitDac_0/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 gnd 2.06fF
C187 9BitDac_0/8BitDac_1/7BitDac_1/V_out7 gnd 2.40fF
C188 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C189 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C190 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C191 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C192 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C193 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C194 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C195 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C196 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C197 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C198 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C199 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C200 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C201 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C202 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C203 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C204 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C205 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C206 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C207 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C208 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C209 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C210 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C211 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C212 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C213 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C214 D0 gnd 203.07fF
C215 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C216 D2 gnd 123.54fF
C217 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C218 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C219 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C220 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C221 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C222 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C223 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C224 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C225 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C226 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C227 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C228 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C229 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C230 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C231 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C232 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C233 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C234 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C235 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C236 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C237 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C238 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C239 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C240 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C241 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C242 9BitDac_0/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 gnd 2.06fF
C243 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C244 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C245 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C246 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C247 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C248 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C249 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C250 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C251 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C252 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C253 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C254 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C255 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C256 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C257 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C258 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C259 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C260 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C261 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C262 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C263 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C264 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C265 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C266 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C267 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C268 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C269 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C270 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C271 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C272 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C273 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C274 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C275 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C276 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C277 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C278 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C279 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C280 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C281 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C282 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C283 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C284 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C285 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C286 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C287 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C288 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C289 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C290 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C291 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C292 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C293 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C294 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C295 9BitDac_1/8BitDac_0/7BitDac_0/6BitDac_1/V_out6 gnd 2.06fF
C296 9BitDac_1/8BitDac_0/7BitDac_1/V_out7 gnd 2.40fF
C297 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C298 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C299 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C300 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C301 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C302 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C303 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C304 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C305 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C306 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C307 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C308 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C309 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C310 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C311 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C312 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C313 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C314 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C315 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C316 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C317 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C318 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C319 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C320 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C321 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C322 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C323 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C324 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C325 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C326 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C327 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C328 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C329 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C330 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C331 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C332 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C333 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C334 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C335 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C336 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C337 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C338 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C339 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C340 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C341 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C342 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C343 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C344 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C345 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C346 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C347 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C348 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C349 9BitDac_1/8BitDac_0/7BitDac_1/6BitDac_1/V_out6 gnd 2.06fF
C350 9BitDac_1/8BitDac_1/V_out8 gnd 2.32fF
C351 9BitDac_1/8BitDac_0/V_out8 gnd 2.04fF
C352 9BitDac_1/8BitDac_1/R_in8 gnd 2.05fF
C353 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C354 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C355 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C356 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C357 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C358 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C359 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C360 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C361 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C362 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C363 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C364 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C365 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C366 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C367 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C368 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C369 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C370 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C371 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C372 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C373 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C374 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C375 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C376 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C377 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C378 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C379 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C380 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C381 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C382 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C383 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C384 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C385 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C386 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C387 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C388 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C389 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C390 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C391 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C392 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C393 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C394 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C395 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C396 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C397 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C398 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C399 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C400 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C401 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C402 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C403 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C404 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C405 9BitDac_1/8BitDac_1/7BitDac_0/6BitDac_1/V_out6 gnd 2.06fF
C406 9BitDac_1/8BitDac_1/7BitDac_1/V_out7 gnd 2.40fF
C407 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C408 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C409 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C410 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C411 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C412 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C413 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C414 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C415 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C416 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C417 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C418 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C419 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C420 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C421 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C422 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C423 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C424 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C425 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C426 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C427 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C428 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C429 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C430 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C431 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C432 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_0/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C433 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C434 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C435 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.35fF
C436 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C437 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/V_out4 gnd 2.39fF
C438 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C439 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C440 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C441 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C442 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C443 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C444 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C445 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_0/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C446 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C447 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/V_out3 gnd 2.43fF
C448 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_0/2BitDac_0/V_out2 gnd 2.39fF
C449 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/V_out3 gnd 2.17fF
C450 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/V_out4 gnd 2.39fF
C451 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C452 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_0/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C453 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_1/V_out2 gnd 2.11fF
C454 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/V_out3 gnd 2.43fF
C455 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_0/2BitDac_0/V_out2 gnd 2.36fF
C456 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/V_out3 gnd 2.17fF
C457 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_1/V_out2 gnd 2.11fF
C458 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/5BitDac_1/4BitDac_1/3BitDac_1/2BitDac_0/V_out2 gnd 2.35fF
C459 9BitDac_1/8BitDac_1/7BitDac_1/6BitDac_1/V_out6 gnd 2.06fF
C460 V_out10 gnd 23.54fF



valpha  R_in10 Gnd 3.3
vbeta  VA Gnd 3.3
vzero D0 Gnd pulse(0 1.8 0.1m 60p 60p 0.1m 0.2m)
vone  D1 Gnd pulse(0 1.8 0.2m 60p 60p 0.2m 0.4m)
vtwo  D2 Gnd pulse(0 1.8 0.4m 60p 60p 0.4m 0.8m)
vthree D3 Gnd pulse(0 1.8 0.8m 60p 60p 0.8m 1.6m)
vfour D4 Gnd pulse (0 1.8 1.6m 60p 60p 1.6m 3.2m)
vfive D5 Gnd pulse (0 1.8 3.2m 60p 60p 3.2m 6.4m)
vsix D6 Gnd pulse (0 1.8 6.4m 60p 60p 6.4m 12.8m)
vseven D7 Gnd pulse (0 1.8 12.8m 60p 60p 12.8m 25.6m)
veight D8 Gnd pulse (0 1.8 25.6m 60p 60p 25.6m 51.2m)
vnine D9 Gnd pulse (0 1.8 51.2m 60p 60p 51.2m 102.4m)
.tran 0.01m 102.4m
.control
run

plot V(V_out10) V(D0)

.endc
.end