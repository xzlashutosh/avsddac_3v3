magic
tech scmos
timestamp 1598795390
<< metal1 >>
rect 331 3297 338 3304
rect 16 3225 21 3227
rect 136 3203 200 3210
rect 331 3177 337 3297
rect 825 3269 831 3276
rect 825 3255 830 3269
rect 825 3248 831 3255
rect 612 3224 1310 3227
rect 481 1573 484 1577
rect 612 1575 616 3224
rect 628 3214 671 3219
rect 604 1572 617 1575
rect 19 -1 23 0
rect 628 -1 632 3214
rect 666 3212 671 3214
rect 1258 1559 1265 1562
rect 1261 1334 1265 1559
rect 1307 1397 1310 3224
rect 1309 1361 1318 1365
rect 1428 1364 1432 1367
rect 1261 1331 1310 1334
rect 19 -5 632 -1
rect 669 -14 673 -13
<< m2contact >>
rect 480 1569 485 1573
rect 1130 1556 1135 1560
rect 1304 1361 1309 1365
<< metal2 >>
rect 481 3245 484 3246
rect 481 3242 1133 3245
rect 481 1573 484 3242
rect 1130 1560 1133 3242
rect 1304 1365 1308 3235
<< m3contact >>
rect 331 3297 338 3304
rect 825 3269 831 3276
rect 825 3248 831 3255
rect 136 3203 143 3210
rect 196 3203 201 3210
rect 331 3177 337 3184
<< metal3 >>
rect 338 3297 987 3304
rect 175 3269 825 3275
rect 40 3218 44 3223
rect 40 3212 61 3218
rect 58 3210 61 3212
rect 58 3204 136 3210
rect 175 3161 179 3269
rect 185 3259 838 3262
rect 185 3162 188 3259
rect 201 3204 694 3210
rect 690 3203 694 3204
rect 331 2455 337 3177
rect 825 3148 829 3248
rect 835 3149 838 3259
rect 981 2441 987 3297
<< metal4 >>
rect 163 3284 821 3288
rect 163 3216 171 3284
rect 813 3203 821 3284
use 6BitDac  6BitDac_0
timestamp 1598764253
transform 1 0 877 0 1 1539
box -877 -1539 -269 1686
use 6BitDac  6BitDac_1
timestamp 1598764253
transform 1 0 1527 0 1 1526
box -877 -1539 -269 1686
use switchNew  switchNew_0
timestamp 1598622215
transform 1 0 1241 0 1 1325
box 69 6 187 75
<< labels >>
rlabel metal1 16 3227 21 3227 5 R_in7
rlabel metal1 1432 1364 1432 1367 7 V_out7
rlabel metal2 1304 3235 1308 3235 5 D6!
rlabel metal1 669 -14 673 -14 1 R_out7
rlabel metal1 333 3244 333 3244 1 D4!
rlabel metal3 40 3218 44 3218 1 D0!
rlabel metal3 40 3223 44 3223 1 D0!
rlabel metal3 185 3262 188 3262 1 D2!
rlabel metal4 163 3288 171 3288 5 D3!
rlabel metal3 175 3275 179 3275 1 D1!
rlabel metal2 481 3246 484 3246 5 D5!
rlabel metal1 828 3264 828 3264 1 D1!
rlabel metal3 835 3262 838 3262 1 D2!
rlabel metal3 331 3177 337 3177 1 D4!
rlabel metal3 344 3304 350 3304 5 D4!
<< end >>
