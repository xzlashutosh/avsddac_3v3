magic
tech scmos
timestamp 1598619523
<< nwell >>
rect 83 -34 141 -7
rect 147 -34 176 -7
rect 180 -69 213 -47
rect 219 -80 278 -53
rect 284 -80 312 -53
rect 80 -125 140 -98
rect 146 -125 174 -98
rect 316 -115 349 -93
rect 178 -160 211 -138
<< ntransistor >>
rect 193 -25 195 -20
rect 96 -54 98 -49
rect 126 -60 128 -55
rect 161 -61 163 -56
rect 329 -71 331 -66
rect 232 -100 234 -95
rect 262 -106 264 -101
rect 297 -107 299 -102
rect 191 -116 193 -111
rect 93 -145 95 -140
rect 123 -151 125 -146
rect 159 -152 161 -147
<< ptransistor >>
rect 96 -28 98 -18
rect 126 -28 128 -18
rect 161 -28 163 -18
rect 193 -63 195 -53
rect 232 -74 234 -64
rect 262 -74 264 -64
rect 297 -74 299 -64
rect 329 -109 331 -99
rect 93 -119 95 -109
rect 123 -119 125 -109
rect 159 -119 161 -109
rect 191 -154 193 -144
<< ndiffusion >>
rect 186 -21 193 -20
rect 186 -25 187 -21
rect 191 -25 193 -21
rect 195 -24 197 -20
rect 201 -24 202 -20
rect 195 -25 202 -24
rect 89 -53 90 -49
rect 94 -53 96 -49
rect 89 -54 96 -53
rect 98 -53 100 -49
rect 104 -53 105 -49
rect 98 -54 105 -53
rect 119 -59 120 -55
rect 124 -59 126 -55
rect 119 -60 126 -59
rect 128 -59 130 -55
rect 134 -59 135 -55
rect 128 -60 135 -59
rect 154 -60 155 -56
rect 159 -60 161 -56
rect 154 -61 161 -60
rect 163 -60 165 -56
rect 169 -60 170 -56
rect 163 -61 170 -60
rect 322 -67 329 -66
rect 322 -71 323 -67
rect 327 -71 329 -67
rect 331 -70 333 -66
rect 337 -70 338 -66
rect 331 -71 338 -70
rect 225 -99 226 -95
rect 230 -99 232 -95
rect 225 -100 232 -99
rect 234 -99 236 -95
rect 240 -99 241 -95
rect 234 -100 241 -99
rect 255 -105 256 -101
rect 260 -105 262 -101
rect 255 -106 262 -105
rect 264 -105 266 -101
rect 270 -105 271 -101
rect 264 -106 271 -105
rect 290 -106 291 -102
rect 295 -106 297 -102
rect 290 -107 297 -106
rect 299 -106 301 -102
rect 305 -106 306 -102
rect 299 -107 306 -106
rect 184 -112 191 -111
rect 184 -116 185 -112
rect 189 -116 191 -112
rect 193 -115 195 -111
rect 199 -115 200 -111
rect 193 -116 200 -115
rect 86 -144 87 -140
rect 91 -144 93 -140
rect 86 -145 93 -144
rect 95 -144 97 -140
rect 101 -144 102 -140
rect 95 -145 102 -144
rect 116 -150 117 -146
rect 121 -150 123 -146
rect 116 -151 123 -150
rect 125 -150 127 -146
rect 131 -150 132 -146
rect 125 -151 132 -150
rect 152 -151 153 -147
rect 157 -151 159 -147
rect 152 -152 159 -151
rect 161 -151 163 -147
rect 167 -151 168 -147
rect 161 -152 168 -151
<< pdiffusion >>
rect 89 -21 96 -18
rect 89 -25 90 -21
rect 94 -25 96 -21
rect 89 -28 96 -25
rect 98 -21 105 -18
rect 98 -25 100 -21
rect 104 -25 105 -21
rect 98 -28 105 -25
rect 119 -21 126 -18
rect 119 -25 120 -21
rect 124 -25 126 -21
rect 119 -28 126 -25
rect 128 -21 135 -18
rect 128 -25 130 -21
rect 134 -25 135 -21
rect 128 -28 135 -25
rect 154 -21 161 -18
rect 154 -25 155 -21
rect 159 -25 161 -21
rect 154 -28 161 -25
rect 163 -21 170 -18
rect 163 -25 165 -21
rect 169 -25 170 -21
rect 163 -28 170 -25
rect 186 -56 193 -53
rect 186 -60 187 -56
rect 191 -60 193 -56
rect 186 -63 193 -60
rect 195 -56 202 -53
rect 195 -60 197 -56
rect 201 -60 202 -56
rect 195 -63 202 -60
rect 225 -67 232 -64
rect 225 -71 226 -67
rect 230 -71 232 -67
rect 225 -74 232 -71
rect 234 -67 241 -64
rect 234 -71 236 -67
rect 240 -71 241 -67
rect 234 -74 241 -71
rect 255 -67 262 -64
rect 255 -71 256 -67
rect 260 -71 262 -67
rect 255 -74 262 -71
rect 264 -67 271 -64
rect 264 -71 266 -67
rect 270 -71 271 -67
rect 264 -74 271 -71
rect 290 -67 297 -64
rect 290 -71 291 -67
rect 295 -71 297 -67
rect 290 -74 297 -71
rect 299 -67 306 -64
rect 299 -71 301 -67
rect 305 -71 306 -67
rect 299 -74 306 -71
rect 322 -102 329 -99
rect 322 -106 323 -102
rect 327 -106 329 -102
rect 322 -109 329 -106
rect 331 -102 338 -99
rect 331 -106 333 -102
rect 337 -106 338 -102
rect 331 -109 338 -106
rect 86 -112 93 -109
rect 86 -116 87 -112
rect 91 -116 93 -112
rect 86 -119 93 -116
rect 95 -112 102 -109
rect 95 -116 97 -112
rect 101 -116 102 -112
rect 95 -119 102 -116
rect 116 -112 123 -109
rect 116 -116 117 -112
rect 121 -116 123 -112
rect 116 -119 123 -116
rect 125 -112 132 -109
rect 125 -116 127 -112
rect 131 -116 132 -112
rect 125 -119 132 -116
rect 152 -112 159 -109
rect 152 -116 153 -112
rect 157 -116 159 -112
rect 152 -119 159 -116
rect 161 -112 168 -109
rect 161 -116 163 -112
rect 167 -116 168 -112
rect 161 -119 168 -116
rect 184 -147 191 -144
rect 184 -151 185 -147
rect 189 -151 191 -147
rect 184 -154 191 -151
rect 193 -147 200 -144
rect 193 -151 195 -147
rect 199 -151 200 -147
rect 193 -154 200 -151
<< ndcontact >>
rect 187 -25 191 -21
rect 197 -24 201 -20
rect 90 -53 94 -49
rect 100 -53 104 -49
rect 120 -59 124 -55
rect 130 -59 134 -55
rect 155 -60 159 -56
rect 165 -60 169 -56
rect 323 -71 327 -67
rect 333 -70 337 -66
rect 226 -99 230 -95
rect 236 -99 240 -95
rect 256 -105 260 -101
rect 266 -105 270 -101
rect 291 -106 295 -102
rect 301 -106 305 -102
rect 185 -116 189 -112
rect 195 -115 199 -111
rect 87 -144 91 -140
rect 97 -144 101 -140
rect 117 -150 121 -146
rect 127 -150 131 -146
rect 153 -151 157 -147
rect 163 -151 167 -147
<< pdcontact >>
rect 90 -25 94 -21
rect 100 -25 104 -21
rect 120 -25 124 -21
rect 130 -25 134 -21
rect 155 -25 159 -21
rect 165 -25 169 -21
rect 187 -60 191 -56
rect 197 -60 201 -56
rect 226 -71 230 -67
rect 236 -71 240 -67
rect 256 -71 260 -67
rect 266 -71 270 -67
rect 291 -71 295 -67
rect 301 -71 305 -67
rect 323 -106 327 -102
rect 333 -106 337 -102
rect 87 -116 91 -112
rect 97 -116 101 -112
rect 117 -116 121 -112
rect 127 -116 131 -112
rect 153 -116 157 -112
rect 163 -116 167 -112
rect 185 -151 189 -147
rect 195 -151 199 -147
<< psubstratepcontact >>
rect 90 -69 94 -65
rect 98 -69 102 -65
rect 120 -69 124 -65
rect 128 -69 132 -65
rect 226 -115 230 -111
rect 234 -115 238 -111
rect 256 -115 260 -111
rect 264 -115 268 -111
rect 87 -160 91 -156
rect 95 -160 99 -156
rect 117 -160 121 -156
rect 125 -160 129 -156
<< nsubstratencontact >>
rect 90 -14 94 -10
rect 98 -14 102 -10
rect 120 -14 124 -10
rect 128 -14 132 -10
rect 155 -14 159 -10
rect 206 -56 210 -52
rect 226 -60 230 -56
rect 234 -60 238 -56
rect 256 -60 260 -56
rect 264 -60 268 -56
rect 291 -60 295 -56
rect 87 -105 91 -101
rect 95 -105 99 -101
rect 103 -105 107 -101
rect 117 -105 121 -101
rect 125 -105 129 -101
rect 153 -105 157 -101
rect 342 -102 346 -98
rect 204 -147 208 -143
<< polysilicon >>
rect 96 -18 98 -16
rect 126 -18 128 -16
rect 161 -18 163 -16
rect 193 -20 195 -18
rect 96 -38 98 -28
rect 97 -42 98 -38
rect 126 -41 128 -28
rect 161 -41 163 -28
rect 193 -33 195 -25
rect 194 -37 195 -33
rect 96 -49 98 -42
rect 127 -45 128 -41
rect 162 -45 163 -41
rect 96 -56 98 -54
rect 126 -55 128 -45
rect 161 -56 163 -45
rect 193 -53 195 -37
rect 126 -62 128 -60
rect 161 -63 163 -61
rect 193 -65 195 -63
rect 232 -64 234 -62
rect 262 -64 264 -62
rect 297 -64 299 -62
rect 329 -66 331 -64
rect 232 -84 234 -74
rect 233 -88 234 -84
rect 262 -87 264 -74
rect 297 -87 299 -74
rect 329 -79 331 -71
rect 330 -83 331 -79
rect 232 -95 234 -88
rect 263 -91 264 -87
rect 298 -91 299 -87
rect 232 -102 234 -100
rect 262 -101 264 -91
rect 297 -102 299 -91
rect 329 -99 331 -83
rect 93 -109 95 -107
rect 123 -109 125 -107
rect 159 -109 161 -107
rect 262 -108 264 -106
rect 297 -109 299 -107
rect 191 -111 193 -109
rect 329 -111 331 -109
rect 93 -129 95 -119
rect 94 -133 95 -129
rect 123 -132 125 -119
rect 159 -132 161 -119
rect 191 -124 193 -116
rect 192 -128 193 -124
rect 93 -140 95 -133
rect 124 -136 125 -132
rect 160 -136 161 -132
rect 93 -147 95 -145
rect 123 -146 125 -136
rect 159 -147 161 -136
rect 191 -144 193 -128
rect 123 -153 125 -151
rect 159 -154 161 -152
rect 191 -156 193 -154
<< polycontact >>
rect 93 -42 97 -38
rect 190 -37 194 -33
rect 123 -45 127 -41
rect 158 -45 162 -41
rect 229 -88 233 -84
rect 326 -83 330 -79
rect 259 -91 263 -87
rect 294 -91 298 -87
rect 90 -133 94 -129
rect 188 -128 192 -124
rect 120 -136 124 -132
rect 156 -136 160 -132
<< metal1 >>
rect 54 15 59 27
rect 71 -2 76 7
rect 53 -3 76 -2
rect 53 -6 154 -3
rect 53 -7 76 -6
rect 53 -33 58 -7
rect 151 -10 154 -6
rect 94 -14 98 -10
rect 102 -14 120 -10
rect 124 -14 128 -10
rect 132 -14 134 -10
rect 151 -14 155 -10
rect 159 -14 201 -10
rect 90 -21 94 -14
rect 120 -21 124 -14
rect 155 -21 159 -14
rect 197 -20 201 -14
rect 70 -72 75 -41
rect 89 -42 93 -38
rect 100 -41 104 -25
rect 130 -34 134 -25
rect 134 -38 150 -34
rect 165 -41 169 -25
rect 187 -27 191 -25
rect 187 -30 201 -27
rect 181 -37 190 -34
rect 181 -38 194 -37
rect 197 -36 201 -30
rect 197 -39 223 -36
rect 197 -41 201 -39
rect 100 -45 123 -41
rect 127 -45 158 -41
rect 165 -45 201 -41
rect 100 -49 104 -45
rect 90 -65 94 -53
rect 130 -55 134 -52
rect 165 -56 169 -45
rect 197 -56 201 -45
rect 206 -52 210 -39
rect 219 -49 223 -39
rect 219 -52 290 -49
rect 287 -56 290 -52
rect 120 -65 124 -59
rect 230 -60 234 -56
rect 238 -60 256 -56
rect 260 -60 264 -56
rect 268 -60 270 -56
rect 287 -60 291 -56
rect 295 -60 337 -56
rect 155 -65 159 -60
rect 187 -65 191 -60
rect 94 -69 98 -65
rect 102 -69 120 -65
rect 124 -69 128 -65
rect 132 -69 133 -65
rect 148 -69 191 -65
rect 226 -67 230 -60
rect 256 -67 260 -60
rect 291 -67 295 -60
rect 333 -66 337 -60
rect 148 -72 151 -69
rect 53 -75 151 -72
rect 53 -82 58 -75
rect 227 -88 229 -84
rect 236 -87 240 -71
rect 266 -80 270 -71
rect 270 -84 286 -80
rect 301 -87 305 -71
rect 323 -73 327 -71
rect 323 -76 337 -73
rect 317 -83 326 -80
rect 317 -84 330 -83
rect 333 -82 337 -76
rect 333 -85 351 -82
rect 333 -87 337 -85
rect 70 -94 75 -90
rect 236 -91 259 -87
rect 263 -91 294 -87
rect 301 -91 337 -87
rect 70 -97 152 -94
rect 236 -95 240 -91
rect 70 -109 74 -97
rect 149 -101 152 -97
rect 53 -113 74 -109
rect 91 -105 95 -101
rect 99 -105 103 -101
rect 107 -105 117 -101
rect 121 -105 125 -101
rect 129 -105 131 -101
rect 149 -105 153 -101
rect 157 -105 199 -101
rect 87 -112 91 -105
rect 117 -112 121 -105
rect 153 -112 157 -105
rect 195 -111 199 -105
rect 53 -132 58 -113
rect 86 -133 90 -129
rect 97 -132 101 -116
rect 127 -125 131 -116
rect 131 -129 148 -125
rect 163 -132 167 -116
rect 226 -111 230 -99
rect 266 -101 270 -98
rect 301 -102 305 -91
rect 333 -102 337 -91
rect 342 -98 346 -85
rect 256 -111 260 -105
rect 291 -111 295 -106
rect 323 -111 327 -106
rect 230 -115 234 -111
rect 238 -115 256 -111
rect 260 -115 264 -111
rect 268 -115 269 -111
rect 284 -115 327 -111
rect 185 -118 189 -116
rect 284 -118 287 -115
rect 185 -121 199 -118
rect 179 -128 188 -125
rect 179 -129 192 -128
rect 195 -127 199 -121
rect 212 -121 287 -118
rect 212 -127 216 -121
rect 195 -130 216 -127
rect 195 -132 199 -130
rect 97 -136 120 -132
rect 124 -136 156 -132
rect 163 -136 199 -132
rect 97 -140 101 -136
rect 70 -163 75 -140
rect 87 -156 91 -144
rect 127 -146 131 -143
rect 163 -147 167 -136
rect 195 -147 199 -136
rect 204 -143 208 -130
rect 117 -156 121 -150
rect 153 -156 157 -151
rect 185 -156 189 -151
rect 91 -160 95 -156
rect 99 -160 117 -156
rect 121 -160 125 -156
rect 129 -160 130 -156
rect 146 -160 189 -156
rect 103 -163 106 -160
rect 146 -163 149 -160
rect 70 -166 149 -163
<< m2contact >>
rect 130 -38 134 -34
rect 150 -38 154 -34
rect 177 -38 181 -34
rect 130 -52 134 -48
rect 266 -84 270 -80
rect 286 -84 290 -80
rect 313 -84 317 -80
rect 266 -98 270 -94
rect 127 -129 131 -125
rect 148 -129 152 -125
rect 175 -129 179 -125
rect 127 -143 131 -139
<< metal2 >>
rect 154 -38 177 -34
rect 130 -48 134 -38
rect 290 -84 313 -80
rect 266 -94 270 -84
rect 152 -129 175 -125
rect 127 -139 131 -129
<< pseudo_rpoly >>
rect 89 -69 90 -65
rect 225 -115 226 -111
rect 86 -160 87 -156
use resistor  resistor_0
timestamp 1598617915
transform 1 0 62 0 1 9
box -9 -7 15 11
use resistor  resistor_1
timestamp 1598617915
transform 1 0 61 0 1 -39
box -9 -7 15 11
use resistor  resistor_2
timestamp 1598617915
transform 1 0 61 0 1 -88
box -9 -7 15 11
use resistor  resistor_3
timestamp 1598617915
transform 1 0 61 0 1 -138
box -9 -7 15 11
<< labels >>
rlabel metal1 262 -113 262 -113 1 gnd!
rlabel metal1 232 -113 232 -113 1 gnd!
rlabel metal1 227 -88 227 -84 1 D1
rlabel metal1 54 27 59 27 4 va
rlabel metal1 74 -4 74 -4 1 alpha
rlabel metal1 73 -73 73 -73 1 beta
rlabel metal1 72 -111 72 -111 1 gamma
rlabel metal1 73 -158 73 -158 1 delta
rlabel metal1 96 -67 96 -67 1 gnd!
rlabel metal1 126 -67 126 -67 1 gnd!
rlabel metal1 89 -42 89 -38 1 D0
rlabel metal1 86 -133 86 -129 1 D0
rlabel metal1 93 -158 93 -158 1 gnd!
rlabel metal1 123 -158 123 -158 1 gnd!
rlabel metal1 351 -85 351 -82 7 V_out
rlabel metal1 106 -10 109 -10 1 Vdd!
rlabel metal1 108 -101 111 -101 1 Vdd!
rlabel metal1 242 -56 245 -56 1 Vdd!
<< end >>
