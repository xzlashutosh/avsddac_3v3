magic
tech scmos
timestamp 1599295951
<< metal1 >>
rect 3022 3366 6005 3369
rect 2363 3359 2999 3360
rect 2339 3356 2999 3359
rect 2334 3279 2338 3337
rect 16 3269 21 3273
rect 3022 1612 3025 3366
rect 3053 3288 3058 3356
rect 3053 3285 3215 3288
rect 3211 3274 3215 3285
rect 3211 3269 3248 3274
rect 3252 3269 3258 3274
rect 3020 1609 3025 1612
rect 3057 3258 3084 3263
rect 3057 31 3061 3258
rect 6002 1822 6005 3366
rect 6002 1819 6025 1822
rect 6027 1783 6033 1787
rect 6143 1786 6147 1789
rect 6023 1740 6026 1756
rect 6023 1737 6083 1740
rect 6080 1603 6083 1737
rect 3056 25 3061 31
rect 3056 1 3060 25
rect 2166 0 3060 1
rect 2162 -3 3060 0
rect 5225 -7 5229 -6
<< m2contact >>
rect 2334 3354 2339 3360
rect 2999 3356 3006 3360
rect 2334 3337 2339 3343
rect 2451 3284 2463 3290
rect 2502 3285 2514 3291
rect 2334 3274 2341 3279
rect 3051 3356 3058 3360
rect 3248 3269 3252 3276
rect 6022 1783 6027 1787
<< metal2 >>
rect 2891 3376 5959 3379
rect 2334 3343 2339 3354
rect 2891 3351 2894 3376
rect 3006 3356 3051 3360
rect 3123 3350 4346 3353
rect 2797 3328 2859 3331
rect 3123 3331 3126 3350
rect 2913 3328 3126 3331
rect 3211 3332 3329 3336
rect 3211 3296 3215 3332
rect 2965 3292 3215 3296
rect 481 3280 484 3285
rect 2463 3285 2502 3290
rect 2463 3284 2507 3285
rect 1304 3269 1309 3272
rect 2626 3257 2750 3260
rect 2965 3260 2968 3292
rect 2918 3257 2968 3260
rect 3325 3263 3329 3332
rect 4343 3325 4346 3350
rect 4400 3325 4418 3326
rect 4343 3323 4418 3325
rect 4343 3322 4420 3323
rect 5860 3322 5864 3362
rect 5956 3349 5959 3376
rect 5954 3346 5959 3349
rect 4400 3321 4420 3322
rect 3544 3274 3547 3279
rect 4367 3263 4372 3266
rect 3325 3259 3547 3263
rect 6022 1787 6025 3220
<< m3contact >>
rect 2859 3328 2867 3332
rect 2905 3328 2913 3332
rect 2334 3274 2341 3279
rect 2750 3257 2755 3262
rect 2913 3257 2918 3262
rect 3248 3269 3252 3276
<< metal3 >>
rect 344 3338 350 3346
rect 3179 3339 3384 3346
rect 2867 3328 2905 3331
rect 3179 3319 3186 3339
rect 3377 3332 3384 3339
rect 3407 3335 3413 3338
rect 3377 3325 3428 3332
rect 2474 3312 3186 3319
rect 175 3309 179 3312
rect 3238 3303 3242 3306
rect 185 3298 188 3300
rect 3248 3293 3251 3294
rect 2502 3290 2514 3291
rect 2318 3284 2463 3290
rect 2502 3286 2945 3290
rect 2502 3285 2514 3286
rect 2328 3274 2334 3277
rect 40 3259 44 3264
rect 2755 3257 2913 3260
rect 2941 3236 2945 3286
rect 3032 3268 3177 3272
rect 3032 3236 3036 3268
rect 3103 3255 3107 3259
rect 3173 3257 3177 3268
rect 3173 3253 3242 3257
rect 2941 3232 3036 3236
rect 2187 3219 2203 3225
rect 3090 68 3094 81
rect 3090 64 3095 68
rect 2170 6 2174 60
rect 3091 6 3095 64
rect 2170 2 3100 6
<< metal4 >>
rect 163 3327 171 3330
rect 3226 3321 3234 3324
rect 2306 3299 3230 3303
<< metal5 >>
rect 2995 3277 3122 3282
rect 115 3223 122 3229
rect 2284 3216 2292 3224
rect 2995 3172 3000 3277
rect 3117 3226 3122 3277
rect 3117 3221 3143 3226
rect 2349 3167 3000 3172
rect 5991 1825 6059 1829
rect 5991 1644 5995 1825
rect 6055 1822 6059 1825
<< metal6 >>
rect 6047 1745 6101 1750
rect 6096 1522 6101 1745
rect 5993 1517 6101 1522
rect 2220 -6 2233 -5
rect 2220 -9 2234 -6
rect 2228 -12 2234 -9
rect 3212 -12 3218 8
rect 2228 -18 3218 -12
rect 5239 -40 5246 -9
use 8BitDac  8BitDac_0
timestamp 1599268620
transform 1 0 0 0 1 20
box 0 -29 3020 3332
use switchNew  switchNew_0
timestamp 1599222484
transform 1 0 5956 0 1 1747
box 69 -1 187 81
use 8BitDac  8BitDac_1
timestamp 1599268620
transform 1 0 3063 0 1 14
box 0 -29 3020 3332
<< labels >>
rlabel metal1 6147 1786 6147 1789 7 V_out9
rlabel metal1 16 3273 21 3273 1 R_in9
rlabel metal2 6022 3214 6025 3214 1 D8!
rlabel metal5 115 3223 122 3223 1 VA
rlabel metal4 163 3330 171 3330 1 D3
rlabel metal3 175 3312 179 3312 1 D1
rlabel metal3 185 3300 188 3300 1 D2
rlabel metal3 344 3346 350 3346 1 D4
rlabel metal2 481 3285 484 3285 1 D5
rlabel metal2 1304 3272 1309 3272 1 D6
rlabel metal3 3103 3259 3107 3259 1 D0
rlabel metal4 3226 3324 3234 3324 1 D3
rlabel metal3 3238 3306 3242 3306 1 D1
rlabel metal3 3248 3294 3251 3294 1 D2
rlabel metal3 3407 3338 3413 3338 1 D4
rlabel metal2 3544 3279 3547 3279 1 D5
rlabel metal2 4367 3266 4372 3266 1 D6
rlabel metal2 5954 3349 5957 3349 1 D7
rlabel metal2 6022 3220 6025 3220 1 D8
rlabel metal5 2284 3224 2292 3224 1 VA
rlabel metal1 5225 -7 5229 -7 1 R_out9
rlabel metal6 5239 -40 5245 -40 1 gnd
rlabel metal3 40 3264 44 3264 1 D0
<< end >>
