magic
tech scmos
timestamp 1599268620
<< metal1 >>
rect 8 799 13 800
rect 169 378 172 382
rect 308 10 311 384
rect 308 7 323 10
rect 308 6 322 7
rect 0 -8 22 0
rect 327 -29 329 -25
rect 439 -26 441 -23
rect 314 -59 330 -56
rect 314 -422 317 -59
rect 162 -428 164 -424
rect 301 -425 317 -422
rect 10 -808 14 -806
<< metal3 >>
rect 32 787 36 790
rect 167 734 171 736
rect 177 734 180 735
rect 159 87 163 88
rect 157 83 165 87
rect 26 -8 29 45
rect 24 -13 29 -8
rect 24 -19 28 -13
rect 159 -72 163 83
rect 172 -12 175 189
rect 171 -15 175 -12
rect 169 -72 174 -15
<< metal5 >>
rect 133 775 141 795
rect 79 84 83 90
rect 79 -10 85 84
rect 209 14 355 19
rect 79 -16 133 -10
rect 125 -31 133 -16
rect 209 -60 214 14
rect 185 -64 214 -60
rect 193 -65 214 -64
<< metal6 >>
rect 33 -119 43 9
rect 343 -68 350 -61
rect 344 -166 350 -68
rect 180 -172 350 -166
use 4BitDac  4BitDac_0
timestamp 1599268620
transform 1 0 10 0 1 395
box -10 -395 301 404
use 4BitDac  4BitDac_1
timestamp 1599268620
transform 1 0 2 0 1 -411
box -10 -395 301 404
use switchNew  switchNew_0
timestamp 1599222484
transform 1 0 252 0 1 -65
box 69 -1 187 81
<< labels >>
rlabel metal1 441 -26 441 -23 7 V_out5
rlabel metal3 167 736 171 736 1 D1!
rlabel metal3 177 735 180 735 1 D2!
rlabel metal1 8 800 13 800 5 R_in5
rlabel metal3 32 790 36 790 1 D0!
rlabel metal1 10 -808 14 -808 1 R_out5
<< end >>
