magic
tech scmos
timestamp 1599268620
<< metal1 >>
rect -861 1685 -856 1686
rect -703 1263 -700 1267
rect -428 859 -416 862
rect -710 457 -707 461
rect -860 68 -855 82
rect -419 69 -416 859
rect -397 104 -393 789
rect -419 66 -390 69
rect -393 30 -382 34
rect -273 33 -269 36
rect -421 0 -389 3
rect -421 -5 -390 0
rect -704 -352 -699 -348
rect -421 -753 -413 -5
rect -427 -756 -413 -753
rect -708 -1158 -706 -1154
rect -858 -1539 -854 -1536
<< m2contact >>
rect -708 1263 -703 1267
rect -555 856 -542 860
rect -721 456 -710 461
rect -711 262 -702 270
rect -397 97 -393 104
rect -397 30 -393 34
rect -711 -352 -704 -348
rect -551 -759 -541 -755
rect -716 -1159 -708 -1154
<< metal2 >>
rect -397 34 -393 97
<< m3contact >>
rect -708 1263 -703 1267
rect -555 856 -542 860
rect -721 456 -710 461
rect -711 262 -702 270
rect -711 -352 -704 -348
rect -551 -759 -541 -755
rect -716 -1159 -708 -1154
<< metal3 >>
rect -837 1681 -833 1682
rect -702 1638 -698 1639
rect -692 1620 -689 1622
rect -555 860 -550 1533
rect -555 844 -551 856
rect -555 840 -545 844
rect -549 398 -545 840
rect -551 394 -545 398
rect -705 270 -702 271
rect -711 260 -702 262
rect -711 253 -708 260
rect -711 250 -665 253
rect -711 245 -708 250
rect -668 213 -665 250
rect -668 210 -663 213
rect -850 70 -847 125
rect -850 66 -832 70
rect -836 63 -832 66
rect -716 24 -712 167
rect -666 30 -663 210
rect -691 27 -663 30
rect -716 20 -697 24
rect -691 5 -688 27
rect -551 -755 -547 394
<< m4contact >>
rect -708 1263 -703 1267
rect -721 456 -710 461
rect -711 -352 -704 -348
rect -716 -1159 -708 -1154
<< metal4 >>
rect -715 1357 -710 1672
rect -715 1352 -703 1357
rect -708 1267 -703 1352
rect -708 1250 -703 1263
rect -716 1245 -703 1250
rect -716 984 -711 1245
rect -726 979 -711 984
rect -726 968 -721 979
rect -726 963 -716 968
rect -721 461 -716 963
rect -721 370 -716 456
rect -725 365 -716 370
rect -725 346 -720 365
rect -725 341 -717 346
rect -722 181 -717 341
rect -731 176 -717 181
rect -731 125 -726 176
rect -731 120 -698 125
rect -703 41 -698 120
rect -710 36 -698 41
rect -710 -38 -705 36
rect -714 -43 -705 -38
rect -714 -63 -709 -43
rect -714 -68 -706 -63
rect -711 -228 -706 -68
rect -722 -233 -706 -228
rect -722 -251 -717 -233
rect -722 -256 -709 -251
rect -714 -267 -709 -256
rect -714 -270 -708 -267
rect -711 -348 -708 -270
rect -704 -352 -699 -348
rect -711 -632 -708 -352
rect -719 -635 -708 -632
rect -719 -673 -716 -635
rect -719 -676 -707 -673
rect -710 -800 -707 -676
rect -716 -803 -707 -800
rect -716 -1154 -713 -803
<< metal5 >>
rect -790 169 -747 174
rect -790 166 -726 169
rect -755 161 -726 166
rect -734 153 -726 161
rect -734 145 -711 153
rect -719 102 -711 145
rect -719 94 -705 102
rect -713 73 -705 94
rect -735 65 -705 73
rect -444 77 -356 85
rect -735 58 -727 65
rect -444 58 -436 77
rect -360 71 -356 77
rect -727 50 -436 58
<< metal6 >>
rect -784 -40 -779 87
rect -827 -43 -816 -40
rect -807 -45 -779 -40
rect -368 -17 -363 -3
rect -368 -90 -362 -17
rect -674 -96 -362 -90
use 5BitDac  5BitDac_0
timestamp 1599268620
transform 1 0 -869 0 1 885
box -8 -808 441 800
use 5BitDac  5BitDac_1
timestamp 1599268620
transform 1 0 -868 0 1 -730
box -8 -808 441 800
use switchNew  switchNew_0
timestamp 1599222484
transform 1 0 -459 0 1 -6
box 69 -1 187 81
<< labels >>
rlabel metal1 -269 33 -269 36 7 V_out6
rlabel metal1 -861 1686 -856 1686 5 R_in6
rlabel metal3 -837 1682 -833 1682 5 D0
rlabel metal3 -702 1639 -698 1639 1 D1
rlabel metal3 -692 1622 -689 1622 1 D2
rlabel metal1 -397 789 -393 789 1 D5
rlabel metal4 -715 1672 -710 1672 1 D3
rlabel metal3 -555 1533 -550 1533 1 D4
rlabel metal1 -858 -1539 -854 -1539 1 R_out6
<< end >>
